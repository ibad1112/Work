magic
tech sky130A
magscale 1 2
timestamp 1606420870
<< nwell >>
rect -1083 -1219 1083 1219
<< pmos >>
rect -887 -1000 -487 1000
rect -429 -1000 -29 1000
rect 29 -1000 429 1000
rect 487 -1000 887 1000
<< pdiff >>
rect -945 988 -887 1000
rect -945 -988 -933 988
rect -899 -988 -887 988
rect -945 -1000 -887 -988
rect -487 988 -429 1000
rect -487 -988 -475 988
rect -441 -988 -429 988
rect -487 -1000 -429 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 429 988 487 1000
rect 429 -988 441 988
rect 475 -988 487 988
rect 429 -1000 487 -988
rect 887 988 945 1000
rect 887 -988 899 988
rect 933 -988 945 988
rect 887 -1000 945 -988
<< pdiffc >>
rect -933 -988 -899 988
rect -475 -988 -441 988
rect -17 -988 17 988
rect 441 -988 475 988
rect 899 -988 933 988
<< nsubdiff >>
rect -1047 1149 -951 1183
rect 951 1149 1047 1183
rect -1047 1087 -1013 1149
rect 1013 1087 1047 1149
rect -1047 -1149 -1013 -1087
rect 1013 -1149 1047 -1087
rect -1047 -1183 -951 -1149
rect 951 -1183 1047 -1149
<< nsubdiffcont >>
rect -951 1149 951 1183
rect -1047 -1087 -1013 1087
rect 1013 -1087 1047 1087
rect -951 -1183 951 -1149
<< poly >>
rect -887 1081 -487 1097
rect -887 1047 -871 1081
rect -503 1047 -487 1081
rect -887 1000 -487 1047
rect -429 1081 -29 1097
rect -429 1047 -413 1081
rect -45 1047 -29 1081
rect -429 1000 -29 1047
rect 29 1081 429 1097
rect 29 1047 45 1081
rect 413 1047 429 1081
rect 29 1000 429 1047
rect 487 1081 887 1097
rect 487 1047 503 1081
rect 871 1047 887 1081
rect 487 1000 887 1047
rect -887 -1047 -487 -1000
rect -887 -1081 -871 -1047
rect -503 -1081 -487 -1047
rect -887 -1097 -487 -1081
rect -429 -1047 -29 -1000
rect -429 -1081 -413 -1047
rect -45 -1081 -29 -1047
rect -429 -1097 -29 -1081
rect 29 -1047 429 -1000
rect 29 -1081 45 -1047
rect 413 -1081 429 -1047
rect 29 -1097 429 -1081
rect 487 -1047 887 -1000
rect 487 -1081 503 -1047
rect 871 -1081 887 -1047
rect 487 -1097 887 -1081
<< polycont >>
rect -871 1047 -503 1081
rect -413 1047 -45 1081
rect 45 1047 413 1081
rect 503 1047 871 1081
rect -871 -1081 -503 -1047
rect -413 -1081 -45 -1047
rect 45 -1081 413 -1047
rect 503 -1081 871 -1047
<< locali >>
rect -1047 1149 -951 1183
rect 951 1149 1047 1183
rect -1047 1087 -1013 1149
rect 1013 1087 1047 1149
rect -887 1047 -871 1081
rect -503 1047 -487 1081
rect -429 1047 -413 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 413 1047 429 1081
rect 487 1047 503 1081
rect 871 1047 887 1081
rect -933 988 -899 1004
rect -933 -1004 -899 -988
rect -475 988 -441 1004
rect -475 -1004 -441 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 441 988 475 1004
rect 441 -1004 475 -988
rect 899 988 933 1004
rect 899 -1004 933 -988
rect -887 -1081 -871 -1047
rect -503 -1081 -487 -1047
rect -429 -1081 -413 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 413 -1081 429 -1047
rect 487 -1081 503 -1047
rect 871 -1081 887 -1047
rect -1047 -1149 -1013 -1087
rect 1013 -1149 1047 -1087
rect -1047 -1183 -951 -1149
rect 951 -1183 1047 -1149
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1030 -1166 1030 1166
string parameters w 10 l 2 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
