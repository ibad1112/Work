magic
tech sky130A
timestamp 1606545195
<< pwell >>
rect -123 -355 123 355
<< nmos >>
rect -25 -250 25 250
<< ndiff >>
rect -54 244 -25 250
rect -54 -244 -48 244
rect -31 -244 -25 244
rect -54 -250 -25 -244
rect 25 244 54 250
rect 25 -244 31 244
rect 48 -244 54 244
rect 25 -250 54 -244
<< ndiffc >>
rect -48 -244 -31 244
rect 31 -244 48 244
<< psubdiff >>
rect -105 320 -57 337
rect 57 320 105 337
rect -105 289 -88 320
rect 88 289 105 320
rect -105 -320 -88 -289
rect 88 -320 105 -289
rect -105 -337 -57 -320
rect 57 -337 105 -320
<< psubdiffcont >>
rect -57 320 57 337
rect -105 -289 -88 289
rect 88 -289 105 289
rect -57 -337 57 -320
<< poly >>
rect -25 286 25 294
rect -25 269 -17 286
rect 17 269 25 286
rect -25 250 25 269
rect -25 -269 25 -250
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -25 -294 25 -286
<< polycont >>
rect -17 269 17 286
rect -17 -286 17 -269
<< locali >>
rect -105 320 -57 337
rect 57 320 105 337
rect -105 289 -88 320
rect 88 289 105 320
rect -25 269 -17 286
rect 17 269 25 286
rect -48 244 -31 252
rect -48 -252 -31 -244
rect 31 244 48 252
rect 31 -252 48 -244
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -105 -320 -88 -289
rect 88 -320 105 -289
rect -105 -337 -57 -320
rect 57 -337 105 -320
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -96 -328 96 328
string parameters w 5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
