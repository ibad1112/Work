magic
tech sky130A
magscale 1 2
timestamp 1606502482
<< nwell >>
rect -396 -261 396 261
<< pmoslvt >>
rect -200 -42 200 42
<< pdiff >>
rect -258 30 -200 42
rect -258 -30 -246 30
rect -212 -30 -200 30
rect -258 -42 -200 -30
rect 200 30 258 42
rect 200 -30 212 30
rect 246 -30 258 30
rect 200 -42 258 -30
<< pdiffc >>
rect -246 -30 -212 30
rect 212 -30 246 30
<< nsubdiff >>
rect -360 191 -264 225
rect 264 191 360 225
rect -360 129 -326 191
rect 326 129 360 191
rect -360 -191 -326 -129
rect 326 -191 360 -129
rect -360 -225 -264 -191
rect 264 -225 360 -191
<< nsubdiffcont >>
rect -264 191 264 225
rect -360 -129 -326 129
rect 326 -129 360 129
rect -264 -225 264 -191
<< poly >>
rect -200 123 200 139
rect -200 89 -184 123
rect 184 89 200 123
rect -200 42 200 89
rect -200 -89 200 -42
rect -200 -123 -184 -89
rect 184 -123 200 -89
rect -200 -139 200 -123
<< polycont >>
rect -184 89 184 123
rect -184 -123 184 -89
<< locali >>
rect -360 191 -264 225
rect 264 191 360 225
rect -360 129 -326 191
rect 326 129 360 191
rect -200 89 -184 123
rect 184 89 200 123
rect -246 30 -212 46
rect -246 -46 -212 -30
rect 212 30 246 46
rect 212 -46 246 -30
rect -200 -123 -184 -89
rect 184 -123 200 -89
rect -360 -191 -326 -129
rect 326 -191 360 -129
rect -360 -225 -264 -191
rect 264 -225 360 -191
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -343 -208 343 208
string parameters w 0.42 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
