magic
tech sky130A
magscale 1 2
timestamp 1606597354
<< nwell >>
rect 15068 3088 18654 3102
rect 15062 2808 18654 3088
rect 15062 2794 18648 2808
<< pwell >>
rect 5358 5118 5894 5146
rect 5284 1898 6636 5118
<< locali >>
rect 7248 2892 7318 2906
rect 7248 2858 7272 2892
rect 7312 2858 7318 2892
rect 7844 2904 7918 2906
rect 7844 2870 7866 2904
rect 7900 2870 7918 2904
rect 7844 2868 7918 2870
rect 7248 2854 7318 2858
rect 12064 2446 12098 2450
rect 12064 2434 12118 2446
rect 12064 2398 12072 2434
rect 12106 2398 12118 2434
rect 12064 2380 12118 2398
rect 12064 2376 12098 2380
<< viali >>
rect 7272 2858 7312 2892
rect 7866 2870 7900 2904
rect 15648 2676 15682 2712
rect 15740 2678 15774 2714
rect 16542 2694 16576 2730
rect 17426 2714 17466 2752
rect 18452 2726 18486 2760
rect 16634 2596 16674 2634
rect 17516 2596 17556 2634
rect 18546 2596 18584 2638
rect 12072 2398 12106 2434
rect 12796 2398 12836 2432
rect 11148 1482 11184 1540
rect 11234 1370 13730 1404
<< metal1 >>
rect 5970 5636 6082 5640
rect 4184 5522 6082 5636
rect 5970 5426 6082 5522
rect 9136 5272 9802 5478
rect 15558 5444 15732 5446
rect 14884 5286 15736 5444
rect 9448 4836 9558 4850
rect 9448 4736 9464 4836
rect 9548 4736 9558 4836
rect 9448 4264 9558 4736
rect 11498 4264 11596 4272
rect 9448 4180 11600 4264
rect 9454 4174 11600 4180
rect 6920 2900 7324 2906
rect 6920 2848 6928 2900
rect 6994 2892 7324 2900
rect 6994 2858 7272 2892
rect 7312 2858 7324 2892
rect 6994 2848 7324 2858
rect 6920 2842 7324 2848
rect 7842 2904 7918 2912
rect 7842 2870 7866 2904
rect 7900 2870 7918 2904
rect 6886 2738 6980 2742
rect 6886 2686 6906 2738
rect 6966 2726 6980 2738
rect 7842 2726 7918 2870
rect 11498 2792 11596 4174
rect 15558 2952 15732 5286
rect 18656 3084 18766 3088
rect 15828 2948 16478 3060
rect 16708 3008 18766 3084
rect 16708 3004 18672 3008
rect 11498 2728 11634 2792
rect 17514 2762 18498 2774
rect 17452 2760 18498 2762
rect 16630 2752 18452 2760
rect 16630 2742 17426 2752
rect 6966 2686 7920 2726
rect 6886 2684 7920 2686
rect 9228 2688 9378 2702
rect 6886 2668 6980 2684
rect 9228 2598 9254 2688
rect 9354 2598 9378 2688
rect 11498 2652 11524 2728
rect 11504 2646 11524 2652
rect 11606 2646 11634 2728
rect 15726 2730 17426 2742
rect 12608 2720 15200 2722
rect 12608 2712 15696 2720
rect 12608 2676 15648 2712
rect 15682 2676 15696 2712
rect 12608 2656 15696 2676
rect 15726 2714 16542 2730
rect 15726 2678 15740 2714
rect 15774 2694 16542 2714
rect 16576 2714 17426 2730
rect 17466 2726 18452 2752
rect 18486 2726 18498 2760
rect 17466 2714 18498 2726
rect 16576 2706 18498 2714
rect 16576 2694 17614 2706
rect 15774 2688 17482 2694
rect 15774 2678 16844 2688
rect 15726 2670 16598 2678
rect 18712 2650 19022 2658
rect 11504 2626 11634 2646
rect 17510 2644 19022 2650
rect 16614 2638 19022 2644
rect 16614 2634 18546 2638
rect 9228 2448 9378 2598
rect 16614 2596 16634 2634
rect 16674 2596 17516 2634
rect 17556 2596 18546 2634
rect 18584 2596 19022 2638
rect 16614 2586 19022 2596
rect 16614 2582 17560 2586
rect 18644 2518 18754 2546
rect 11792 2448 12114 2452
rect 12980 2448 13090 2450
rect 9222 2434 12114 2448
rect 9222 2398 12072 2434
rect 12106 2398 12114 2434
rect 9222 2378 12114 2398
rect 12790 2432 13090 2448
rect 12790 2398 12796 2432
rect 12836 2398 13090 2432
rect 12790 2378 13090 2398
rect 9222 2376 11806 2378
rect 4478 1930 4582 2352
rect 12980 2126 13090 2378
rect 12980 2072 13002 2126
rect 13058 2072 13090 2126
rect 12980 2042 13090 2072
rect 4478 1788 6132 1930
rect 7562 1606 7714 1652
rect 7562 1494 7580 1606
rect 7692 1566 7714 1606
rect 7692 1540 11208 1566
rect 7692 1494 11148 1540
rect 7562 1482 11148 1494
rect 11184 1482 11208 1540
rect 7562 1474 11208 1482
rect 7562 1470 7714 1474
rect 11218 1404 13744 1416
rect 11218 1370 11234 1404
rect 13730 1370 13744 1404
rect 11218 1292 13744 1370
rect 15576 1322 15670 2436
rect 15834 2406 16484 2518
rect 16696 2466 18754 2518
rect 16696 2438 18660 2466
rect 14068 1194 15670 1322
rect 15576 1182 15670 1194
<< via1 >>
rect 7930 4726 8014 4826
rect 9464 4736 9548 4836
rect 7242 4556 7336 4680
rect 7096 2966 7148 3028
rect 7746 2968 7806 3048
rect 8110 2960 8162 3042
rect 6928 2848 6994 2900
rect 6906 2686 6966 2738
rect 9254 2598 9354 2688
rect 11524 2646 11606 2728
rect 7580 2064 7692 2176
rect 13002 2072 13058 2126
rect 9004 1818 9090 1896
rect 7580 1494 7692 1606
rect 10978 1186 11064 1264
<< metal2 >>
rect 7224 4680 7362 5002
rect 7888 4836 9560 4850
rect 7888 4826 9464 4836
rect 7888 4726 7930 4826
rect 8014 4736 9464 4826
rect 9548 4736 9560 4836
rect 8014 4726 9560 4736
rect 7888 4710 9560 4726
rect 7224 4556 7242 4680
rect 7336 4556 7362 4680
rect 5558 3582 5662 3584
rect 1942 3474 3596 3548
rect 1942 3414 3350 3474
rect 3302 3326 3350 3414
rect 3540 3436 3596 3474
rect 3540 3326 3598 3436
rect 5122 3434 5662 3582
rect 3302 3290 3598 3326
rect 5558 3170 5662 3434
rect 7224 3254 7362 4556
rect 6860 3170 6986 3172
rect 5558 3142 6986 3170
rect 5558 3080 6886 3142
rect 6956 3080 6986 3142
rect 5558 3060 6986 3080
rect 6860 3058 6986 3060
rect 7066 3044 7170 3064
rect 7066 2952 7090 3044
rect 7158 2952 7170 3044
rect 4154 2934 4284 2944
rect 7066 2940 7170 2952
rect 4154 2930 7010 2934
rect 4154 2836 4164 2930
rect 4258 2900 7010 2930
rect 4258 2848 6928 2900
rect 6994 2848 7010 2900
rect 4258 2836 7010 2848
rect 4154 2824 7010 2836
rect 4158 2818 7010 2824
rect 6882 2740 6980 2748
rect 6882 2676 6896 2740
rect 6970 2676 6980 2740
rect 6882 2668 6980 2676
rect 7216 2702 7362 3254
rect 8078 3060 8188 3066
rect 7704 3048 8192 3060
rect 7704 3044 7746 3048
rect 7806 3044 8192 3048
rect 7704 2964 7732 3044
rect 7812 3042 8192 3044
rect 7812 2964 8110 3042
rect 7704 2960 8110 2964
rect 8162 2960 8192 3042
rect 7704 2950 8192 2960
rect 11500 2728 11624 2754
rect 7216 2688 9386 2702
rect 7216 2598 9254 2688
rect 9354 2598 9386 2688
rect 7216 2578 9386 2598
rect 7322 2576 9386 2578
rect 11500 2646 11524 2728
rect 11606 2646 11624 2728
rect 7562 2176 7716 2200
rect 7562 2064 7580 2176
rect 7692 2064 7716 2176
rect 7562 1606 7716 2064
rect 11500 2140 11624 2646
rect 12594 2140 13090 2142
rect 11500 2126 13090 2140
rect 11500 2072 13002 2126
rect 13058 2072 13090 2126
rect 11500 2036 13090 2072
rect 7562 1494 7580 1606
rect 7692 1494 7716 1606
rect 7562 1474 7716 1494
rect 8958 1896 9124 1918
rect 8958 1818 9004 1896
rect 9090 1818 9124 1896
rect 8958 1292 9124 1818
rect 8958 1264 11118 1292
rect 8958 1186 10978 1264
rect 11064 1186 11118 1264
rect 8958 1144 11118 1186
<< via2 >>
rect 3350 3326 3540 3474
rect 6886 3080 6956 3142
rect 7090 3028 7158 3044
rect 7090 2966 7096 3028
rect 7096 2966 7148 3028
rect 7148 2966 7158 3028
rect 7090 2952 7158 2966
rect 4164 2836 4258 2930
rect 6896 2738 6970 2740
rect 6896 2686 6906 2738
rect 6906 2686 6966 2738
rect 6966 2686 6970 2738
rect 6896 2676 6970 2686
rect 7732 2968 7746 3044
rect 7746 2968 7806 3044
rect 7806 2968 7812 3044
rect 7732 2964 7812 2968
<< metal3 >>
rect 3274 3474 3634 3554
rect 3274 3326 3350 3474
rect 3540 3326 3634 3474
rect 3274 3302 3634 3326
rect 6866 3142 6988 3170
rect 6866 3080 6886 3142
rect 6956 3080 6988 3142
rect 4066 2930 4290 2960
rect 4066 2836 4164 2930
rect 4258 2836 4290 2930
rect 4066 2806 4290 2836
rect 6866 2740 6988 3080
rect 7100 3066 7892 3068
rect 7064 3044 7892 3066
rect 7064 2952 7090 3044
rect 7158 2964 7732 3044
rect 7812 2964 7892 3044
rect 7158 2952 7892 2964
rect 7064 2938 7186 2952
rect 6866 2676 6896 2740
rect 6970 2676 6988 2740
rect 6866 2656 6988 2676
<< via3 >>
rect 3350 3326 3540 3474
rect 4164 2836 4258 2930
<< metal4 >>
rect 3296 3490 3620 3548
rect 3296 3330 3312 3490
rect 3600 3330 3620 3490
rect 4278 2840 4288 2962
rect 4066 2836 4164 2840
rect 4258 2836 4288 2840
rect 4066 2804 4288 2836
<< via4 >>
rect 3312 3474 3600 3490
rect 3312 3326 3350 3474
rect 3350 3326 3540 3474
rect 3540 3326 3600 3474
rect 3312 3242 3600 3326
rect 3990 2930 4278 3088
rect 3990 2840 4164 2930
rect 4164 2840 4258 2930
rect 4258 2840 4278 2930
<< metal5 >>
rect 3276 3490 3638 3552
rect 3276 3242 3312 3490
rect 3600 3242 3638 3490
rect 3276 3130 3638 3242
rect 3276 3088 4302 3130
rect 3276 2840 3990 3088
rect 4278 2840 4302 3088
rect 3276 2796 4302 2840
rect 3276 2792 3850 2796
use LVDSBias  LVDSBias_0
timestamp 1606277081
transform 1 0 2998 0 1 5224
box -3498 -5224 2404 652
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1606261606
transform 1 0 18380 0 1 2510
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1606261606
transform 1 0 17354 0 1 2492
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1606261606
transform 1 0 16464 0 1 2476
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1606261606
transform 1 0 15566 0 1 2458
box -38 -48 314 592
use LVDS2  LVDS2_0
timestamp 1606076054
transform 1 0 9778 0 1 2844
box -152 -1748 5398 2676
use LVDS1  LVDS1_0
timestamp 1606079819
transform 1 0 5879 0 1 3380
box -53 -1584 3506 2114
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1606272999
transform 1 0 18732 0 1 2508
box -38 -48 130 592
<< labels >>
rlabel metal1 18748 2594 18786 2636 1 OUT
port 1 n
<< end >>
