magic
tech sky130A
magscale 1 2
timestamp 1606607067
<< nwell >>
rect 7862 2528 11846 2532
rect 4870 2486 6072 2490
rect 7862 2486 14424 2528
rect 4870 2238 14424 2486
rect 4870 2218 11846 2238
rect 2628 2202 11846 2218
rect 2628 946 6072 2202
rect 7862 1442 11846 2202
rect 2628 796 4906 946
rect 2544 794 4906 796
rect 524 766 4906 794
rect 524 528 3050 766
rect 524 400 2766 528
rect 524 198 2566 400
rect 524 -10 1014 198
rect 1588 -6 2566 198
rect 6044 78 7972 568
rect 524 -26 900 -10
<< pwell >>
rect 542 -718 1092 -296
rect 1554 -716 2182 -284
rect 2568 -710 3732 -270
rect 4126 -754 4548 -262
rect 7076 -758 7730 -252
<< psubdiff >>
rect 10518 -856 13588 -842
rect 7216 -858 13588 -856
rect 4424 -860 13588 -858
rect -162 -862 762 -860
rect 2590 -862 13588 -860
rect -162 -872 10694 -862
rect -162 -876 5620 -872
rect -162 -880 2944 -876
rect -162 -926 -60 -880
rect -12 -926 98 -880
rect 146 -926 262 -880
rect 310 -926 414 -880
rect 462 -882 774 -880
rect 462 -926 552 -882
rect -162 -928 552 -926
rect 600 -928 774 -882
rect 824 -882 1618 -880
rect 824 -884 1052 -882
rect 824 -928 910 -884
rect -162 -932 910 -928
rect 960 -930 1052 -884
rect 1102 -884 1332 -882
rect 1102 -930 1196 -884
rect 960 -932 1196 -930
rect 1246 -930 1332 -884
rect 1382 -886 1618 -882
rect 1382 -930 1464 -886
rect 1246 -932 1464 -930
rect -162 -934 1464 -932
rect 1514 -928 1618 -886
rect 1668 -882 2598 -880
rect 1668 -886 1968 -882
rect 1668 -928 1794 -886
rect 1514 -934 1794 -928
rect 1848 -930 1968 -886
rect 2022 -884 2598 -882
rect 2022 -886 2254 -884
rect 2022 -930 2116 -886
rect 1848 -934 2116 -930
rect 2170 -932 2254 -886
rect 2308 -888 2598 -884
rect 2308 -932 2414 -888
rect 2170 -934 2414 -932
rect -162 -936 2414 -934
rect 2468 -934 2598 -888
rect 2656 -882 2944 -880
rect 2656 -930 2766 -882
rect 2818 -924 2944 -882
rect 2996 -880 4314 -876
rect 2996 -924 3116 -880
rect 2818 -928 3116 -924
rect 3168 -928 3300 -880
rect 3352 -882 3818 -880
rect 3352 -928 3456 -882
rect 2818 -930 3456 -928
rect 3508 -930 3632 -882
rect 3684 -928 3818 -882
rect 3870 -928 3974 -880
rect 4026 -928 4146 -880
rect 4198 -924 4314 -880
rect 4366 -924 4446 -876
rect 4498 -880 4840 -876
rect 4498 -882 4710 -880
rect 4498 -924 4576 -882
rect 4198 -928 4576 -924
rect 3684 -930 4576 -928
rect 4628 -928 4710 -882
rect 4762 -924 4840 -880
rect 4892 -880 5126 -876
rect 4892 -924 4988 -880
rect 4762 -928 4988 -924
rect 5040 -924 5126 -880
rect 5178 -880 5452 -876
rect 5178 -924 5288 -880
rect 5040 -928 5288 -924
rect 5340 -924 5452 -880
rect 5504 -920 5620 -876
rect 5672 -876 5912 -872
rect 5672 -920 5764 -876
rect 5504 -924 5764 -920
rect 5816 -920 5912 -876
rect 5964 -876 6500 -872
rect 5964 -920 6068 -876
rect 5816 -924 6068 -920
rect 6120 -924 6214 -876
rect 6266 -924 6360 -876
rect 6412 -920 6500 -876
rect 6552 -880 6898 -872
rect 6552 -920 6644 -880
rect 6412 -924 6644 -920
rect 5340 -928 6644 -924
rect 6696 -928 6778 -880
rect 6830 -920 6898 -880
rect 6950 -876 10532 -872
rect 6950 -920 7030 -876
rect 6830 -924 7030 -920
rect 7082 -924 7162 -876
rect 7214 -878 8220 -876
rect 7214 -924 7304 -878
rect 6830 -926 7304 -924
rect 7356 -882 7782 -878
rect 7356 -926 7452 -882
rect 6830 -928 7452 -926
rect 4628 -930 7452 -928
rect 7504 -886 7782 -882
rect 7504 -930 7614 -886
rect 2656 -934 7614 -930
rect 7666 -926 7782 -886
rect 7834 -926 7930 -878
rect 7982 -926 8072 -878
rect 8124 -924 8220 -878
rect 8272 -878 8642 -876
rect 8272 -924 8372 -878
rect 8124 -926 8372 -924
rect 8424 -926 8502 -878
rect 8554 -924 8642 -878
rect 8694 -878 9690 -876
rect 8694 -924 8830 -878
rect 8554 -926 8830 -924
rect 8882 -926 9010 -878
rect 9062 -926 9178 -878
rect 9230 -882 9534 -878
rect 9230 -926 9372 -882
rect 7666 -930 9372 -926
rect 9424 -926 9534 -882
rect 9586 -924 9690 -878
rect 9742 -924 9848 -876
rect 9900 -878 10532 -876
rect 9900 -924 10032 -878
rect 9586 -926 10032 -924
rect 10084 -926 10216 -878
rect 10268 -926 10380 -878
rect 10432 -926 10532 -878
rect 9424 -930 10532 -926
rect 7666 -934 10532 -930
rect 2468 -936 10532 -934
rect 10592 -926 10694 -872
rect 10754 -926 10888 -862
rect 10948 -866 11288 -862
rect 10948 -926 11078 -866
rect 10592 -930 11078 -926
rect 11138 -926 11288 -866
rect 11348 -866 11854 -862
rect 11348 -926 11482 -866
rect 11138 -930 11482 -926
rect 11542 -872 11854 -866
rect 11542 -930 11668 -872
rect 10592 -936 11668 -930
rect 11728 -926 11854 -872
rect 11914 -866 12618 -862
rect 11914 -872 12208 -866
rect 11914 -926 12034 -872
rect 11728 -936 12034 -926
rect 12094 -930 12208 -872
rect 12268 -930 12418 -866
rect 12478 -926 12618 -866
rect 12678 -926 12818 -862
rect 12878 -926 13052 -862
rect 13112 -866 13588 -862
rect 13112 -926 13310 -866
rect 12478 -930 13310 -926
rect 13370 -930 13588 -866
rect 12094 -936 13588 -930
rect -162 -942 13588 -936
rect 1798 -944 13588 -942
rect 1798 -946 2622 -944
rect 4424 -946 13588 -944
rect 7216 -948 9712 -946
rect 10518 -954 13588 -946
<< nsubdiff >>
rect 11790 2442 14300 2448
rect 11746 2436 14300 2442
rect 8046 2426 14300 2436
rect 5736 2418 14300 2426
rect 5736 2414 9522 2418
rect 5736 2412 8396 2414
rect 5736 2410 6864 2412
rect 5736 2366 5848 2410
rect 5900 2406 6290 2410
rect 5900 2366 5996 2406
rect 5736 2362 5996 2366
rect 6048 2362 6124 2406
rect 6176 2366 6290 2406
rect 6342 2408 6864 2410
rect 6342 2366 6428 2408
rect 6176 2364 6428 2366
rect 6480 2406 6716 2408
rect 6480 2364 6578 2406
rect 6176 2362 6578 2364
rect 6630 2364 6716 2406
rect 6768 2368 6864 2408
rect 6916 2410 8396 2412
rect 6916 2408 7284 2410
rect 6916 2406 7148 2408
rect 6916 2368 7002 2406
rect 6768 2364 7002 2368
rect 6630 2362 7002 2364
rect 7054 2364 7148 2406
rect 7200 2366 7284 2408
rect 7336 2408 7550 2410
rect 7336 2366 7412 2408
rect 7200 2364 7412 2366
rect 7464 2366 7550 2408
rect 7602 2366 7682 2410
rect 7734 2408 8396 2410
rect 7734 2406 7982 2408
rect 7734 2366 7822 2406
rect 7464 2364 7822 2366
rect 7054 2362 7822 2364
rect 7874 2364 7982 2406
rect 8034 2364 8134 2408
rect 8186 2364 8270 2408
rect 8322 2370 8396 2408
rect 8448 2370 8560 2414
rect 8612 2412 8828 2414
rect 8612 2370 8704 2412
rect 8322 2368 8704 2370
rect 8756 2370 8828 2412
rect 8880 2370 8992 2414
rect 9044 2412 9318 2414
rect 9044 2370 9150 2412
rect 8756 2368 9150 2370
rect 9202 2370 9318 2412
rect 9370 2374 9522 2414
rect 9574 2374 9676 2418
rect 9728 2374 9850 2418
rect 9902 2374 10050 2418
rect 10102 2374 10200 2418
rect 10252 2374 10364 2418
rect 10416 2374 10514 2418
rect 10566 2414 10860 2418
rect 10566 2374 10652 2414
rect 9370 2370 10652 2374
rect 10704 2374 10860 2414
rect 10912 2374 11008 2418
rect 11060 2412 11452 2418
rect 11060 2374 11220 2412
rect 10704 2370 11220 2374
rect 9202 2368 11220 2370
rect 11272 2374 11452 2412
rect 11504 2414 14300 2418
rect 11504 2374 11636 2414
rect 11272 2370 11636 2374
rect 11688 2372 11818 2414
rect 14232 2372 14300 2414
rect 11688 2370 14300 2372
rect 11272 2368 14300 2370
rect 8322 2364 14300 2368
rect 7874 2362 14300 2364
rect 5736 2350 14300 2362
rect 5736 2344 8054 2350
rect 11746 2348 14300 2350
rect 11746 2346 11986 2348
rect 2700 2144 4864 2166
rect 2700 2140 4024 2144
rect 2700 2134 3124 2140
rect 2700 2082 2810 2134
rect 2862 2082 2960 2134
rect 3012 2088 3124 2134
rect 3176 2138 4024 2140
rect 3176 2134 3728 2138
rect 3176 2088 3284 2134
rect 3012 2082 3284 2088
rect 3336 2082 3440 2134
rect 3492 2082 3582 2134
rect 3634 2086 3728 2134
rect 3780 2086 3866 2138
rect 3918 2092 4024 2138
rect 4076 2140 4864 2144
rect 4076 2092 4174 2140
rect 3918 2088 4174 2092
rect 4226 2088 4346 2140
rect 4398 2088 4502 2140
rect 4554 2088 4684 2140
rect 4736 2088 4864 2140
rect 3918 2086 4864 2088
rect 3634 2082 4864 2086
rect 2700 2058 4864 2082
rect 700 610 770 612
rect 1694 610 2720 612
rect 700 600 2720 610
rect 700 598 1938 600
rect 700 596 1694 598
rect 700 558 742 596
rect 788 558 858 596
rect 904 558 980 596
rect 1026 558 1100 596
rect 1146 558 1216 596
rect 1262 592 1446 596
rect 1262 558 1320 592
rect 700 554 1320 558
rect 1366 558 1446 592
rect 1492 558 1564 596
rect 1610 560 1694 596
rect 1742 596 1938 598
rect 1742 560 1810 596
rect 1610 558 1810 560
rect 1858 562 1938 596
rect 1986 598 2444 600
rect 1986 596 2182 598
rect 1986 562 2068 596
rect 1858 558 2068 562
rect 2116 560 2182 596
rect 2230 560 2306 598
rect 2354 562 2444 598
rect 2492 562 2570 600
rect 2618 562 2720 600
rect 2354 560 2720 562
rect 2116 558 2720 560
rect 1366 554 2720 558
rect 700 546 2720 554
rect 700 540 770 546
rect 1694 544 2720 546
<< psubdiffcont >>
rect -60 -926 -12 -880
rect 98 -926 146 -880
rect 262 -926 310 -880
rect 414 -926 462 -880
rect 552 -928 600 -882
rect 774 -928 824 -880
rect 910 -932 960 -884
rect 1052 -930 1102 -882
rect 1196 -932 1246 -884
rect 1332 -930 1382 -882
rect 1464 -934 1514 -886
rect 1618 -928 1668 -880
rect 1794 -934 1848 -886
rect 1968 -930 2022 -882
rect 2116 -934 2170 -886
rect 2254 -932 2308 -884
rect 2414 -936 2468 -888
rect 2598 -934 2656 -880
rect 2766 -930 2818 -882
rect 2944 -924 2996 -876
rect 3116 -928 3168 -880
rect 3300 -928 3352 -880
rect 3456 -930 3508 -882
rect 3632 -930 3684 -882
rect 3818 -928 3870 -880
rect 3974 -928 4026 -880
rect 4146 -928 4198 -880
rect 4314 -924 4366 -876
rect 4446 -924 4498 -876
rect 4576 -930 4628 -882
rect 4710 -928 4762 -880
rect 4840 -924 4892 -876
rect 4988 -928 5040 -880
rect 5126 -924 5178 -876
rect 5288 -928 5340 -880
rect 5452 -924 5504 -876
rect 5620 -920 5672 -872
rect 5764 -924 5816 -876
rect 5912 -920 5964 -872
rect 6068 -924 6120 -876
rect 6214 -924 6266 -876
rect 6360 -924 6412 -876
rect 6500 -920 6552 -872
rect 6644 -928 6696 -880
rect 6778 -928 6830 -880
rect 6898 -920 6950 -872
rect 7030 -924 7082 -876
rect 7162 -924 7214 -876
rect 7304 -926 7356 -878
rect 7452 -930 7504 -882
rect 7614 -934 7666 -886
rect 7782 -926 7834 -878
rect 7930 -926 7982 -878
rect 8072 -926 8124 -878
rect 8220 -924 8272 -876
rect 8372 -926 8424 -878
rect 8502 -926 8554 -878
rect 8642 -924 8694 -876
rect 8830 -926 8882 -878
rect 9010 -926 9062 -878
rect 9178 -926 9230 -878
rect 9372 -930 9424 -882
rect 9534 -926 9586 -878
rect 9690 -924 9742 -876
rect 9848 -924 9900 -876
rect 10032 -926 10084 -878
rect 10216 -926 10268 -878
rect 10380 -926 10432 -878
rect 10532 -936 10592 -872
rect 10694 -926 10754 -862
rect 10888 -926 10948 -862
rect 11078 -930 11138 -866
rect 11288 -926 11348 -862
rect 11482 -930 11542 -866
rect 11668 -936 11728 -872
rect 11854 -926 11914 -862
rect 12034 -936 12094 -872
rect 12208 -930 12268 -866
rect 12418 -930 12478 -866
rect 12618 -926 12678 -862
rect 12818 -926 12878 -862
rect 13052 -926 13112 -862
rect 13310 -930 13370 -866
<< nsubdiffcont >>
rect 5848 2366 5900 2410
rect 5996 2362 6048 2406
rect 6124 2362 6176 2406
rect 6290 2366 6342 2410
rect 6428 2364 6480 2408
rect 6578 2362 6630 2406
rect 6716 2364 6768 2408
rect 6864 2368 6916 2412
rect 7002 2362 7054 2406
rect 7148 2364 7200 2408
rect 7284 2366 7336 2410
rect 7412 2364 7464 2408
rect 7550 2366 7602 2410
rect 7682 2366 7734 2410
rect 7822 2362 7874 2406
rect 7982 2364 8034 2408
rect 8134 2364 8186 2408
rect 8270 2364 8322 2408
rect 8396 2370 8448 2414
rect 8560 2370 8612 2414
rect 8704 2368 8756 2412
rect 8828 2370 8880 2414
rect 8992 2370 9044 2414
rect 9150 2368 9202 2412
rect 9318 2370 9370 2414
rect 9522 2374 9574 2418
rect 9676 2374 9728 2418
rect 9850 2374 9902 2418
rect 10050 2374 10102 2418
rect 10200 2374 10252 2418
rect 10364 2374 10416 2418
rect 10514 2374 10566 2418
rect 10652 2370 10704 2414
rect 10860 2374 10912 2418
rect 11008 2374 11060 2418
rect 11220 2368 11272 2412
rect 11452 2374 11504 2418
rect 11636 2370 11688 2414
rect 11818 2372 14232 2414
rect 2810 2082 2862 2134
rect 2960 2082 3012 2134
rect 3124 2088 3176 2140
rect 3284 2082 3336 2134
rect 3440 2082 3492 2134
rect 3582 2082 3634 2134
rect 3728 2086 3780 2138
rect 3866 2086 3918 2138
rect 4024 2092 4076 2144
rect 4174 2088 4226 2140
rect 4346 2088 4398 2140
rect 4502 2088 4554 2140
rect 4684 2088 4736 2140
rect 742 558 788 596
rect 858 558 904 596
rect 980 558 1026 596
rect 1100 558 1146 596
rect 1216 558 1262 596
rect 1320 554 1366 592
rect 1446 558 1492 596
rect 1564 558 1610 596
rect 1694 560 1742 598
rect 1810 558 1858 596
rect 1938 562 1986 600
rect 2068 558 2116 596
rect 2182 560 2230 598
rect 2306 560 2354 598
rect 2444 562 2492 600
rect 2570 562 2618 600
<< locali >>
rect 8846 2418 9412 2420
rect 8022 2414 8320 2416
rect 5764 2412 6650 2414
rect 5764 2410 6210 2412
rect 5764 2406 5848 2410
rect 5764 2362 5788 2406
rect 5840 2366 5848 2406
rect 5900 2366 5918 2410
rect 5970 2406 6062 2410
rect 5970 2366 5996 2406
rect 5840 2362 5996 2366
rect 6048 2366 6062 2406
rect 6114 2406 6210 2410
rect 6114 2366 6124 2406
rect 6048 2362 6124 2366
rect 6176 2368 6210 2406
rect 6262 2410 6354 2412
rect 6262 2368 6290 2410
rect 6176 2366 6290 2368
rect 6342 2368 6354 2410
rect 6406 2410 6650 2412
rect 6406 2408 6494 2410
rect 6406 2368 6428 2408
rect 6342 2366 6428 2368
rect 6176 2364 6428 2366
rect 6480 2366 6494 2408
rect 6546 2406 6650 2410
rect 6546 2366 6578 2406
rect 6480 2364 6578 2366
rect 6176 2362 6578 2364
rect 6630 2370 6650 2406
rect 6702 2412 6938 2414
rect 6702 2410 6864 2412
rect 6702 2408 6790 2410
rect 6702 2370 6716 2408
rect 6630 2364 6716 2370
rect 6768 2366 6790 2408
rect 6842 2368 6864 2410
rect 6916 2370 6938 2412
rect 6990 2412 8056 2414
rect 6990 2410 7348 2412
rect 6990 2406 7076 2410
rect 6990 2370 7002 2406
rect 6916 2368 7002 2370
rect 6842 2366 7002 2368
rect 6768 2364 7002 2366
rect 6630 2362 7002 2364
rect 7054 2366 7076 2406
rect 7128 2408 7206 2410
rect 7128 2366 7148 2408
rect 7054 2364 7148 2366
rect 7200 2366 7206 2408
rect 7258 2366 7284 2410
rect 7336 2368 7348 2410
rect 7400 2408 7476 2412
rect 7400 2368 7412 2408
rect 7336 2366 7412 2368
rect 7200 2364 7412 2366
rect 7464 2368 7476 2408
rect 7528 2410 7904 2412
rect 7528 2368 7550 2410
rect 7464 2366 7550 2368
rect 7602 2366 7614 2410
rect 7666 2366 7682 2410
rect 7734 2408 7904 2410
rect 7734 2366 7746 2408
rect 7464 2364 7746 2366
rect 7798 2406 7904 2408
rect 7798 2364 7822 2406
rect 7054 2362 7822 2364
rect 7874 2368 7904 2406
rect 7956 2408 8056 2412
rect 7956 2368 7982 2408
rect 7874 2364 7982 2368
rect 8034 2370 8056 2408
rect 8108 2412 8320 2414
rect 8108 2408 8206 2412
rect 8108 2370 8134 2408
rect 8034 2364 8134 2370
rect 8186 2368 8206 2408
rect 8258 2408 8320 2412
rect 8846 2416 9216 2418
rect 8372 2414 9216 2416
rect 8258 2368 8270 2408
rect 8372 2374 8396 2414
rect 8186 2364 8270 2368
rect 8322 2370 8396 2374
rect 8448 2370 8470 2414
rect 8522 2370 8560 2414
rect 8612 2370 8614 2414
rect 8666 2412 8754 2414
rect 8666 2370 8704 2412
rect 8806 2370 8828 2414
rect 8880 2370 8898 2414
rect 8950 2370 8992 2414
rect 9044 2370 9056 2414
rect 9108 2412 9216 2414
rect 9108 2370 9150 2412
rect 8322 2368 8704 2370
rect 8756 2368 9150 2370
rect 9202 2374 9216 2412
rect 9268 2414 9412 2418
rect 9268 2374 9318 2414
rect 9202 2370 9318 2374
rect 9370 2382 9412 2414
rect 9464 2418 9600 2420
rect 9464 2382 9522 2418
rect 9370 2374 9522 2382
rect 9574 2384 9600 2418
rect 9652 2418 9764 2420
rect 9652 2384 9676 2418
rect 9574 2374 9676 2384
rect 9728 2378 9764 2418
rect 9816 2418 9942 2420
rect 9816 2378 9850 2418
rect 9728 2374 9850 2378
rect 9902 2378 9942 2418
rect 9994 2418 10110 2420
rect 9994 2378 10050 2418
rect 9902 2374 10050 2378
rect 10102 2382 10110 2418
rect 10162 2418 10278 2420
rect 10162 2382 10200 2418
rect 10102 2374 10200 2382
rect 10252 2382 10278 2418
rect 10330 2418 10442 2420
rect 10330 2382 10364 2418
rect 10252 2374 10364 2382
rect 10416 2384 10442 2418
rect 10494 2418 10578 2420
rect 10494 2384 10514 2418
rect 10416 2374 10514 2384
rect 10566 2382 10578 2418
rect 10630 2414 10760 2420
rect 10630 2382 10652 2414
rect 10566 2374 10652 2382
rect 9370 2370 10652 2374
rect 10704 2382 10760 2414
rect 10812 2418 11124 2420
rect 10812 2382 10860 2418
rect 10704 2374 10860 2382
rect 10912 2412 11008 2418
rect 10704 2370 10912 2374
rect 9202 2368 10912 2370
rect 10964 2374 11008 2412
rect 11060 2388 11124 2418
rect 11176 2412 11348 2420
rect 11176 2388 11220 2412
rect 11060 2374 11220 2388
rect 10964 2368 11220 2374
rect 11272 2392 11348 2412
rect 11400 2418 11538 2420
rect 11400 2392 11452 2418
rect 11272 2374 11452 2392
rect 11504 2392 11538 2418
rect 11590 2414 11716 2420
rect 11590 2392 11636 2414
rect 11504 2374 11636 2392
rect 11272 2370 11636 2374
rect 11688 2378 11716 2414
rect 11768 2414 14266 2422
rect 11768 2378 11818 2414
rect 11688 2372 11818 2378
rect 14232 2372 14266 2414
rect 11688 2370 14266 2372
rect 11272 2368 14266 2370
rect 8322 2364 11304 2368
rect 7874 2362 8032 2364
rect 2722 2144 4842 2150
rect 2722 2140 4024 2144
rect 2722 2138 2876 2140
rect 2722 2086 2742 2138
rect 2794 2134 2876 2138
rect 2794 2086 2810 2134
rect 2722 2082 2810 2086
rect 2862 2088 2876 2134
rect 2928 2138 3124 2140
rect 2928 2134 3036 2138
rect 2928 2088 2960 2134
rect 2862 2082 2960 2088
rect 3012 2086 3036 2134
rect 3088 2088 3124 2138
rect 3176 2088 3210 2140
rect 3262 2138 3510 2140
rect 3262 2134 3358 2138
rect 3262 2088 3284 2134
rect 3088 2086 3284 2088
rect 3012 2082 3284 2086
rect 3336 2086 3358 2134
rect 3410 2134 3510 2138
rect 3410 2086 3440 2134
rect 3336 2082 3440 2086
rect 3492 2088 3510 2134
rect 3562 2138 3782 2140
rect 3562 2134 3646 2138
rect 3562 2088 3582 2134
rect 3492 2082 3582 2088
rect 3634 2086 3646 2134
rect 3698 2086 3728 2138
rect 3780 2088 3782 2138
rect 3834 2138 4024 2140
rect 3834 2088 3866 2138
rect 3780 2086 3866 2088
rect 3918 2086 3934 2138
rect 3986 2092 4024 2138
rect 4076 2140 4260 2144
rect 4076 2092 4092 2140
rect 3986 2088 4092 2092
rect 4144 2088 4174 2140
rect 4226 2092 4260 2140
rect 4312 2140 4842 2144
rect 4312 2092 4346 2140
rect 4226 2088 4346 2092
rect 4398 2088 4418 2140
rect 4470 2088 4502 2140
rect 4554 2138 4684 2140
rect 4554 2088 4594 2138
rect 3986 2086 4594 2088
rect 4646 2088 4684 2138
rect 4736 2088 4756 2140
rect 4808 2088 4842 2140
rect 4646 2086 4842 2088
rect 3634 2082 4842 2086
rect 2722 2078 4842 2082
rect 9376 2032 9418 2046
rect 6102 2010 6142 2022
rect 6102 1042 6110 2010
rect 9376 1664 9384 2032
rect 9376 1644 9418 1664
rect 6102 1026 6142 1042
rect 11160 672 13162 682
rect 11160 638 11172 672
rect 13148 638 13162 672
rect 11160 624 13162 638
rect 11058 604 11114 618
rect 704 598 1268 600
rect 704 596 794 598
rect 704 558 742 596
rect 788 560 794 596
rect 840 596 1036 598
rect 840 560 858 596
rect 788 558 858 560
rect 904 594 980 596
rect 904 558 916 594
rect 704 556 916 558
rect 962 558 980 594
rect 1026 560 1036 596
rect 1082 596 1268 598
rect 1082 560 1100 596
rect 1026 558 1100 560
rect 1146 594 1216 596
rect 1146 558 1158 594
rect 962 556 1158 558
rect 1204 558 1216 594
rect 1262 562 1268 596
rect 1314 598 1938 600
rect 1314 596 1694 598
rect 1314 592 1378 596
rect 1314 562 1320 592
rect 1262 558 1320 562
rect 1204 556 1320 558
rect 704 554 1320 556
rect 1366 558 1378 592
rect 1424 558 1446 596
rect 1492 558 1500 596
rect 1546 558 1564 596
rect 1610 558 1632 596
rect 1678 560 1694 596
rect 1742 560 1750 598
rect 1798 596 1874 598
rect 1798 560 1810 596
rect 1678 558 1810 560
rect 1858 560 1874 596
rect 1922 562 1938 598
rect 1986 598 2116 600
rect 1986 562 2000 598
rect 1922 560 2000 562
rect 2048 596 2116 598
rect 2048 560 2068 596
rect 1858 558 2068 560
rect 2164 598 2244 600
rect 2164 562 2182 598
rect 2116 560 2182 562
rect 2230 564 2244 598
rect 2292 598 2444 600
rect 2292 564 2306 598
rect 2230 560 2306 564
rect 2354 596 2444 598
rect 2354 560 2376 596
rect 2116 558 2376 560
rect 2424 562 2444 596
rect 2492 562 2514 600
rect 2562 562 2570 600
rect 2618 596 2710 600
rect 2424 558 2616 562
rect 2664 558 2710 596
rect 11058 570 11062 604
rect 11096 570 11114 604
rect 1366 554 1702 558
rect 704 552 766 554
rect 11058 548 11114 570
rect 204 -492 248 -474
rect 3038 -474 3082 -456
rect 204 -526 208 -492
rect 242 -526 248 -492
rect 3038 -508 3044 -474
rect 3078 -508 3082 -474
rect 5748 -476 5790 -460
rect 204 -546 248 -526
rect 3038 -526 3082 -508
rect 5776 -544 5790 -476
rect 5748 -560 5790 -544
rect 5830 -476 5872 -462
rect 5830 -544 5838 -476
rect 5830 -562 5872 -544
rect 10470 -866 10694 -862
rect 2584 -878 2690 -876
rect 742 -880 2690 -878
rect -144 -882 -60 -880
rect -144 -928 -130 -882
rect -82 -926 -60 -882
rect -12 -882 98 -880
rect -12 -926 20 -882
rect -82 -928 20 -926
rect 68 -926 98 -882
rect 146 -926 178 -880
rect 226 -926 262 -880
rect 310 -882 414 -880
rect 310 -926 326 -882
rect 68 -928 326 -926
rect 374 -926 414 -882
rect 462 -882 710 -880
rect 462 -926 476 -882
rect 374 -928 476 -926
rect 524 -928 552 -882
rect 600 -928 622 -882
rect 670 -928 710 -882
rect 756 -928 774 -880
rect 824 -884 976 -880
rect 824 -928 838 -884
rect -144 -932 838 -928
rect 888 -932 910 -884
rect 960 -928 976 -884
rect 1026 -882 1548 -880
rect 1026 -928 1052 -882
rect 960 -930 1052 -928
rect 1102 -930 1118 -882
rect 1168 -884 1332 -882
rect 1168 -930 1196 -884
rect 960 -932 1196 -930
rect 1246 -886 1332 -884
rect 1246 -932 1260 -886
rect 742 -934 1260 -932
rect 1310 -930 1332 -886
rect 1382 -930 1406 -882
rect 1456 -886 1548 -882
rect 1456 -930 1464 -886
rect 1310 -934 1464 -930
rect 1514 -928 1548 -886
rect 1598 -928 1618 -880
rect 1668 -928 1720 -880
rect 1770 -882 2598 -880
rect 1770 -884 1968 -882
rect 1770 -886 1886 -884
rect 1770 -928 1794 -886
rect 1514 -934 1794 -928
rect 1848 -932 1886 -886
rect 1940 -930 1968 -884
rect 2022 -930 2040 -882
rect 2094 -886 2188 -882
rect 2094 -930 2116 -886
rect 1940 -932 2116 -930
rect 1848 -934 2116 -932
rect 2170 -930 2188 -886
rect 2242 -884 2330 -882
rect 2242 -930 2254 -884
rect 2170 -932 2254 -930
rect 2308 -930 2330 -884
rect 2384 -888 2500 -882
rect 2384 -930 2414 -888
rect 2308 -932 2414 -930
rect 2170 -934 2414 -932
rect 742 -936 2414 -934
rect 2468 -930 2500 -888
rect 2554 -930 2598 -882
rect 2468 -934 2598 -930
rect 2656 -928 2690 -880
rect 2748 -882 2858 -876
rect 2748 -928 2766 -882
rect 2656 -930 2766 -928
rect 2818 -928 2858 -882
rect 2916 -924 2944 -876
rect 2996 -924 3030 -876
rect 2916 -928 3030 -924
rect 3088 -880 3208 -876
rect 3088 -928 3116 -880
rect 3168 -928 3208 -880
rect 3266 -880 3380 -876
rect 3266 -928 3300 -880
rect 3352 -928 3380 -880
rect 2818 -930 3380 -928
rect 3438 -880 3730 -876
rect 3438 -882 3546 -880
rect 3438 -930 3456 -882
rect 3508 -930 3546 -882
rect 2656 -934 3546 -930
rect 3604 -882 3730 -880
rect 3604 -930 3632 -882
rect 3684 -930 3730 -882
rect 3788 -880 3900 -876
rect 3788 -928 3818 -880
rect 3870 -928 3900 -880
rect 3788 -930 3900 -928
rect 3958 -880 4060 -876
rect 3958 -928 3974 -880
rect 4026 -928 4060 -880
rect 4118 -880 4240 -876
rect 4118 -928 4146 -880
rect 4198 -928 4240 -880
rect 4402 -876 4638 -872
rect 4298 -924 4314 -876
rect 4366 -924 4384 -876
rect 4436 -924 4446 -876
rect 4498 -924 4508 -876
rect 4560 -882 4638 -876
rect 4560 -924 4576 -882
rect 4298 -928 4576 -924
rect 3958 -930 4576 -928
rect 4628 -918 4638 -882
rect 4690 -880 4776 -872
rect 4690 -918 4710 -880
rect 4628 -928 4710 -918
rect 4762 -918 4776 -880
rect 4828 -876 4912 -872
rect 4828 -918 4840 -876
rect 4762 -924 4840 -918
rect 4892 -918 4912 -876
rect 4964 -880 5054 -872
rect 4964 -918 4988 -880
rect 4892 -924 4988 -918
rect 4762 -928 4988 -924
rect 5040 -918 5054 -880
rect 5106 -876 5542 -872
rect 5106 -918 5126 -876
rect 5040 -924 5126 -918
rect 5178 -924 5212 -876
rect 5264 -880 5380 -876
rect 5264 -924 5288 -880
rect 5040 -928 5288 -924
rect 5340 -924 5380 -880
rect 5432 -924 5452 -876
rect 5504 -918 5542 -876
rect 5594 -918 5620 -872
rect 5504 -920 5620 -918
rect 5672 -876 5836 -872
rect 5672 -920 5682 -876
rect 5504 -924 5682 -920
rect 5734 -924 5764 -876
rect 5816 -920 5836 -876
rect 5888 -920 5912 -872
rect 5964 -918 5992 -872
rect 7650 -872 9262 -870
rect 10470 -872 10606 -866
rect 6044 -876 6284 -872
rect 6044 -918 6068 -876
rect 5964 -920 6068 -918
rect 5816 -924 6068 -920
rect 6120 -924 6142 -876
rect 6194 -924 6214 -876
rect 6266 -920 6284 -876
rect 6336 -876 6432 -872
rect 6336 -920 6360 -876
rect 6266 -924 6360 -920
rect 6412 -920 6432 -876
rect 6484 -920 6500 -872
rect 6552 -876 6898 -872
rect 6552 -920 6576 -876
rect 6412 -924 6576 -920
rect 6628 -880 6710 -876
rect 6628 -924 6644 -880
rect 5340 -928 6644 -924
rect 6696 -924 6710 -880
rect 6762 -880 6898 -876
rect 6762 -924 6778 -880
rect 6696 -928 6778 -924
rect 6830 -882 6898 -880
rect 6830 -928 6840 -882
rect 4628 -930 6840 -928
rect 6892 -920 6898 -882
rect 6950 -874 9262 -872
rect 6950 -876 10454 -874
rect 6950 -882 7030 -876
rect 6950 -920 6958 -882
rect 6892 -930 6958 -920
rect 7010 -924 7030 -882
rect 7082 -882 7162 -876
rect 7082 -924 7092 -882
rect 7010 -930 7092 -924
rect 7144 -924 7162 -882
rect 7214 -878 7532 -876
rect 7214 -924 7230 -878
rect 7144 -926 7230 -924
rect 7282 -926 7304 -878
rect 7356 -926 7376 -878
rect 7428 -882 7532 -878
rect 7428 -926 7452 -882
rect 7144 -930 7452 -926
rect 7504 -924 7532 -882
rect 7584 -886 7702 -876
rect 7584 -924 7614 -886
rect 7504 -930 7614 -924
rect 3604 -932 7614 -930
rect 3604 -934 4410 -932
rect 6056 -934 7614 -932
rect 7666 -924 7702 -886
rect 7754 -878 7998 -876
rect 7754 -924 7782 -878
rect 7666 -926 7782 -924
rect 7834 -880 7930 -878
rect 7834 -926 7860 -880
rect 7666 -928 7860 -926
rect 7912 -926 7930 -880
rect 7982 -924 7998 -878
rect 8050 -878 8220 -876
rect 8050 -924 8072 -878
rect 7982 -926 8072 -924
rect 8124 -926 8142 -878
rect 8194 -924 8220 -878
rect 8272 -878 8642 -876
rect 8272 -880 8372 -878
rect 8272 -924 8298 -880
rect 8194 -926 8298 -924
rect 7912 -928 8298 -926
rect 8350 -926 8372 -880
rect 8424 -880 8502 -878
rect 8424 -926 8434 -880
rect 8350 -928 8434 -926
rect 8486 -926 8502 -880
rect 8554 -880 8642 -878
rect 8554 -926 8576 -880
rect 8486 -928 8576 -926
rect 8628 -924 8642 -880
rect 8694 -878 9264 -876
rect 8694 -886 8830 -878
rect 8694 -924 8724 -886
rect 8628 -928 8724 -924
rect 7666 -934 8724 -928
rect 8776 -926 8830 -886
rect 8882 -880 9010 -878
rect 8882 -926 8928 -880
rect 8776 -928 8928 -926
rect 8980 -926 9010 -880
rect 9062 -886 9178 -878
rect 9062 -926 9100 -886
rect 8980 -928 9100 -926
rect 8776 -934 9100 -928
rect 9152 -926 9178 -886
rect 9230 -924 9264 -878
rect 9316 -882 9462 -876
rect 9316 -924 9372 -882
rect 9230 -926 9372 -924
rect 9152 -930 9372 -926
rect 9424 -924 9462 -882
rect 9514 -878 9690 -876
rect 9514 -924 9534 -878
rect 9424 -926 9534 -924
rect 9586 -880 9690 -878
rect 9586 -926 9630 -880
rect 9424 -928 9630 -926
rect 9682 -924 9690 -880
rect 9742 -878 9848 -876
rect 9742 -924 9768 -878
rect 9682 -926 9768 -924
rect 9820 -924 9848 -878
rect 9900 -924 9934 -876
rect 9986 -878 10454 -876
rect 9986 -924 10032 -878
rect 9820 -926 10032 -924
rect 10084 -926 10128 -878
rect 10180 -926 10216 -878
rect 10268 -882 10380 -878
rect 10268 -926 10290 -882
rect 9682 -928 10290 -926
rect 9424 -930 10290 -928
rect 10342 -926 10380 -882
rect 10432 -926 10454 -878
rect 10342 -930 10454 -926
rect 9152 -934 10454 -930
rect 2468 -936 2592 -934
rect 10514 -936 10532 -872
rect 10592 -930 10606 -872
rect 10666 -926 10694 -866
rect 10754 -926 10790 -862
rect 10850 -926 10888 -862
rect 10948 -926 11000 -862
rect 11060 -866 11196 -862
rect 11060 -926 11078 -866
rect 10666 -930 11078 -926
rect 11138 -926 11196 -866
rect 11256 -926 11288 -862
rect 11348 -926 11386 -862
rect 11446 -866 11586 -862
rect 11446 -926 11482 -866
rect 11138 -930 11482 -926
rect 11542 -920 11586 -866
rect 11646 -866 11854 -862
rect 11646 -872 11770 -866
rect 11646 -920 11668 -872
rect 11542 -930 11668 -920
rect 10592 -936 11668 -930
rect 11728 -930 11770 -872
rect 11830 -926 11854 -866
rect 11914 -926 11946 -862
rect 12006 -866 12618 -862
rect 12006 -872 12208 -866
rect 12006 -926 12034 -872
rect 11830 -930 12034 -926
rect 11728 -936 12034 -930
rect 12094 -936 12116 -872
rect 12176 -930 12208 -872
rect 12268 -930 12330 -866
rect 12390 -930 12418 -866
rect 12478 -930 12526 -866
rect 12586 -926 12618 -866
rect 12678 -876 12818 -862
rect 12678 -926 12710 -876
rect 12586 -930 12710 -926
rect 12176 -936 12710 -930
rect 12770 -926 12818 -876
rect 12878 -926 12950 -862
rect 13010 -926 13052 -862
rect 13112 -866 13432 -862
rect 13112 -926 13174 -866
rect 12770 -930 13174 -926
rect 13234 -930 13310 -866
rect 13370 -926 13432 -866
rect 13492 -926 13554 -862
rect 13370 -930 13554 -926
rect 12770 -936 13554 -930
<< viali >>
rect 5788 2362 5840 2406
rect 5918 2366 5970 2410
rect 6062 2366 6114 2410
rect 6210 2368 6262 2412
rect 6354 2368 6406 2412
rect 6494 2366 6546 2410
rect 6650 2370 6702 2414
rect 6790 2366 6842 2410
rect 6938 2370 6990 2414
rect 7076 2366 7128 2410
rect 7206 2366 7258 2410
rect 7348 2368 7400 2412
rect 7476 2368 7528 2412
rect 7614 2366 7666 2410
rect 7746 2364 7798 2408
rect 7904 2368 7956 2412
rect 8056 2370 8108 2414
rect 8206 2368 8258 2412
rect 8320 2408 8372 2418
rect 8320 2374 8322 2408
rect 8322 2374 8372 2408
rect 8470 2370 8522 2414
rect 8614 2370 8666 2414
rect 8754 2412 8806 2414
rect 8754 2370 8756 2412
rect 8756 2370 8806 2412
rect 8898 2370 8950 2414
rect 9056 2370 9108 2414
rect 9216 2374 9268 2418
rect 9412 2382 9464 2426
rect 9600 2384 9652 2428
rect 9764 2378 9816 2422
rect 9942 2378 9994 2422
rect 10110 2382 10162 2426
rect 10278 2382 10330 2426
rect 10442 2384 10494 2428
rect 10578 2382 10630 2426
rect 10760 2382 10812 2426
rect 10912 2368 10964 2412
rect 11124 2388 11176 2432
rect 11348 2392 11400 2436
rect 11538 2392 11590 2436
rect 11716 2378 11768 2422
rect 11818 2372 14232 2414
rect 6122 2150 7796 2184
rect 9402 2172 11576 2206
rect 11976 2170 14150 2204
rect 2742 2086 2794 2138
rect 2876 2088 2928 2140
rect 3036 2086 3088 2138
rect 3210 2088 3262 2140
rect 3358 2086 3410 2138
rect 3510 2088 3562 2140
rect 3646 2086 3698 2138
rect 3782 2088 3834 2140
rect 3934 2086 3986 2138
rect 4092 2088 4144 2140
rect 4260 2092 4312 2144
rect 4418 2088 4470 2140
rect 4594 2086 4646 2138
rect 4756 2088 4808 2140
rect 6221 2036 7697 2070
rect 9501 2058 11477 2092
rect 12075 2056 14051 2090
rect 3002 1866 4676 1900
rect 3101 1752 4577 1786
rect 3008 756 3042 1724
rect 4636 756 4670 1724
rect 6110 1042 6144 2010
rect 9384 1664 9418 2032
rect 14110 1660 14144 2028
rect 9501 1600 11477 1634
rect 12075 1598 14051 1632
rect 6221 978 7697 1012
rect 3101 694 4577 728
rect 11172 638 13148 672
rect 794 560 840 598
rect 916 556 962 594
rect 1036 560 1082 598
rect 1158 556 1204 594
rect 1268 562 1314 600
rect 1378 558 1424 596
rect 1500 558 1546 596
rect 1632 558 1678 596
rect 1750 560 1798 598
rect 1874 560 1922 598
rect 2000 560 2048 598
rect 2116 562 2164 600
rect 2244 564 2292 602
rect 2376 558 2424 596
rect 2514 562 2562 600
rect 2616 562 2618 596
rect 2618 562 2664 596
rect 2616 558 2664 562
rect 11062 570 11096 604
rect 5568 484 5942 518
rect 8020 498 8394 532
rect 11174 524 13150 558
rect 1132 344 1506 378
rect 5667 370 5843 404
rect 8119 384 8295 418
rect 11084 410 13240 444
rect 2102 336 2476 370
rect 5902 304 5936 342
rect 8354 318 8388 356
rect 1231 230 1407 264
rect 2201 222 2377 256
rect 1138 186 1172 220
rect 3498 216 3558 250
rect 5667 242 5843 276
rect 8119 256 8295 290
rect 2108 178 2142 212
rect 1231 142 1407 176
rect 3414 172 3448 206
rect 2201 134 2377 168
rect 3498 128 3558 162
rect 3408 14 3648 48
rect 11030 -142 13406 -108
rect 306 -482 366 -448
rect 1282 -474 1388 -440
rect 2262 -470 2368 -436
rect 3142 -464 3202 -430
rect 3932 -456 3992 -422
rect 4710 -448 5686 -414
rect 5928 -448 6904 -414
rect 7828 -446 8804 -412
rect 9046 -446 10022 -412
rect 208 -526 242 -492
rect 1198 -518 1232 -484
rect 2178 -514 2212 -480
rect 3044 -508 3078 -474
rect 3838 -498 3872 -464
rect 306 -570 366 -536
rect 1282 -562 1388 -528
rect 2262 -558 2368 -524
rect 3142 -552 3202 -518
rect 3932 -544 3992 -510
rect 5742 -544 5776 -476
rect 5838 -544 5872 -476
rect 6954 -544 6988 -476
rect 7744 -542 7778 -474
rect 8854 -542 8888 -474
rect 8962 -542 8996 -474
rect 10946 -538 10980 -170
rect 4710 -606 5686 -572
rect 5928 -606 6904 -572
rect 7828 -604 8804 -570
rect 9046 -604 10022 -570
rect 11030 -600 13406 -566
rect 216 -684 456 -650
rect 1192 -676 1478 -642
rect 2172 -672 2458 -638
rect 3052 -666 3292 -632
rect 3842 -658 4082 -624
rect 4620 -720 6994 -686
rect 7738 -718 10112 -684
rect 10940 -714 13496 -680
rect -130 -928 -82 -882
rect 20 -928 68 -882
rect 178 -926 226 -880
rect 326 -928 374 -882
rect 476 -928 524 -882
rect 622 -928 670 -882
rect 710 -928 756 -880
rect 838 -932 888 -884
rect 976 -928 1026 -880
rect 1118 -930 1168 -882
rect 1260 -934 1310 -886
rect 1406 -930 1456 -882
rect 1548 -928 1598 -880
rect 1720 -928 1770 -880
rect 1886 -932 1940 -884
rect 2040 -930 2094 -882
rect 2188 -930 2242 -882
rect 2330 -930 2384 -882
rect 2500 -930 2554 -882
rect 2690 -928 2748 -874
rect 2858 -928 2916 -874
rect 3030 -928 3088 -874
rect 3208 -928 3266 -874
rect 3380 -930 3438 -876
rect 3546 -934 3604 -880
rect 3730 -930 3788 -876
rect 3900 -930 3958 -876
rect 4060 -928 4118 -874
rect 4240 -928 4298 -874
rect 4384 -924 4436 -876
rect 4508 -924 4560 -876
rect 4638 -918 4690 -870
rect 4776 -918 4828 -870
rect 4912 -918 4964 -870
rect 5054 -918 5106 -870
rect 5212 -924 5264 -876
rect 5380 -924 5432 -876
rect 5542 -918 5594 -870
rect 5682 -924 5734 -876
rect 5836 -920 5888 -872
rect 5992 -918 6044 -870
rect 6142 -924 6194 -876
rect 6284 -920 6336 -872
rect 6432 -920 6484 -872
rect 6576 -924 6628 -876
rect 6710 -924 6762 -876
rect 6840 -930 6892 -882
rect 6958 -930 7010 -882
rect 7092 -930 7144 -882
rect 7230 -926 7282 -878
rect 7376 -926 7428 -878
rect 7532 -924 7584 -876
rect 7702 -924 7754 -876
rect 7860 -928 7912 -880
rect 7998 -924 8050 -876
rect 8142 -926 8194 -878
rect 8298 -928 8350 -880
rect 8434 -928 8486 -880
rect 8576 -928 8628 -880
rect 8724 -934 8776 -886
rect 8928 -928 8980 -880
rect 9100 -934 9152 -886
rect 9264 -924 9316 -876
rect 9462 -924 9514 -876
rect 9630 -928 9682 -880
rect 9768 -926 9820 -878
rect 9934 -924 9986 -876
rect 10128 -926 10180 -878
rect 10290 -930 10342 -882
rect 10454 -936 10514 -872
rect 10606 -930 10666 -866
rect 10790 -926 10850 -862
rect 11000 -926 11060 -862
rect 11196 -926 11256 -862
rect 11386 -926 11446 -862
rect 11586 -920 11646 -856
rect 11770 -930 11830 -866
rect 11946 -926 12006 -862
rect 12116 -936 12176 -872
rect 12330 -930 12390 -866
rect 12526 -930 12586 -866
rect 12710 -940 12770 -876
rect 12950 -926 13010 -862
rect 13174 -930 13234 -866
rect 13432 -926 13492 -862
<< metal1 >>
rect 11856 2474 14386 2476
rect 9040 2470 14386 2474
rect 5700 2466 8116 2468
rect 4866 2464 8116 2466
rect 8834 2464 14386 2470
rect 4866 2436 14386 2464
rect 4866 2432 11348 2436
rect 4866 2428 11124 2432
rect 4866 2426 9600 2428
rect 4866 2418 9412 2426
rect 4866 2414 8320 2418
rect 4866 2412 6650 2414
rect 4866 2410 6210 2412
rect 4866 2406 5918 2410
rect 4866 2362 5788 2406
rect 5840 2366 5918 2406
rect 5970 2366 6062 2410
rect 6114 2368 6210 2410
rect 6262 2368 6354 2412
rect 6406 2410 6650 2412
rect 6406 2368 6494 2410
rect 6114 2366 6494 2368
rect 6546 2370 6650 2410
rect 6702 2410 6938 2414
rect 6702 2370 6790 2410
rect 6546 2366 6790 2370
rect 6842 2370 6938 2410
rect 6990 2412 8056 2414
rect 6990 2410 7348 2412
rect 6990 2370 7076 2410
rect 6842 2366 7076 2370
rect 7128 2366 7206 2410
rect 7258 2368 7348 2410
rect 7400 2368 7476 2412
rect 7528 2410 7904 2412
rect 7528 2368 7614 2410
rect 7258 2366 7614 2368
rect 7666 2408 7904 2410
rect 7666 2366 7746 2408
rect 5840 2364 7746 2366
rect 7798 2368 7904 2408
rect 7956 2370 8056 2412
rect 8108 2412 8320 2414
rect 8108 2370 8206 2412
rect 7956 2368 8206 2370
rect 8258 2374 8320 2412
rect 8372 2414 9216 2418
rect 8372 2374 8470 2414
rect 8258 2370 8470 2374
rect 8522 2370 8614 2414
rect 8666 2370 8754 2414
rect 8806 2370 8898 2414
rect 8950 2370 9056 2414
rect 9108 2374 9216 2414
rect 9268 2382 9412 2418
rect 9464 2384 9600 2426
rect 9652 2426 10442 2428
rect 9652 2422 10110 2426
rect 9652 2384 9764 2422
rect 9464 2382 9764 2384
rect 9268 2378 9764 2382
rect 9816 2378 9942 2422
rect 9994 2382 10110 2422
rect 10162 2382 10278 2426
rect 10330 2384 10442 2426
rect 10494 2426 11124 2428
rect 10494 2384 10578 2426
rect 10330 2382 10578 2384
rect 10630 2382 10760 2426
rect 10812 2412 11124 2426
rect 10812 2382 10912 2412
rect 9994 2378 10912 2382
rect 9268 2374 10912 2378
rect 9108 2370 10912 2374
rect 8258 2368 10912 2370
rect 10964 2388 11124 2412
rect 11176 2392 11348 2432
rect 11400 2392 11538 2436
rect 11590 2422 14386 2436
rect 11590 2392 11716 2422
rect 11176 2388 11716 2392
rect 10964 2378 11716 2388
rect 11768 2414 14386 2422
rect 11768 2378 11818 2414
rect 10964 2372 11818 2378
rect 14232 2372 14386 2414
rect 10964 2368 14386 2372
rect 7798 2364 14386 2368
rect 5840 2362 14386 2364
rect 4866 2312 14386 2362
rect 4866 2308 8116 2312
rect 8834 2310 14386 2312
rect 8834 2308 9144 2310
rect 4866 2188 5734 2308
rect 2684 2186 5734 2188
rect 2668 2168 5734 2186
rect 6100 2184 7810 2308
rect 2668 2144 4898 2168
rect 2668 2140 4260 2144
rect 2668 2138 2876 2140
rect 2668 2086 2742 2138
rect 2794 2088 2876 2138
rect 2928 2138 3210 2140
rect 2928 2088 3036 2138
rect 2794 2086 3036 2088
rect 3088 2088 3210 2138
rect 3262 2138 3510 2140
rect 3262 2088 3358 2138
rect 3088 2086 3358 2088
rect 3410 2088 3510 2138
rect 3562 2138 3782 2140
rect 3562 2088 3646 2138
rect 3410 2086 3646 2088
rect 3698 2088 3782 2138
rect 3834 2138 4092 2140
rect 3834 2088 3934 2138
rect 3698 2086 3934 2088
rect 3986 2088 4092 2138
rect 4144 2092 4260 2140
rect 4312 2140 4898 2144
rect 4312 2092 4418 2140
rect 4144 2088 4418 2092
rect 4470 2138 4756 2140
rect 4470 2088 4594 2138
rect 3986 2086 4594 2088
rect 4646 2088 4756 2138
rect 4808 2088 4898 2140
rect 6100 2150 6122 2184
rect 7796 2150 7810 2184
rect 6100 2138 7810 2150
rect 6206 2088 7714 2138
rect 4646 2086 4898 2088
rect 2668 2026 4898 2086
rect 6210 2070 7714 2088
rect 6210 2036 6221 2070
rect 7697 2036 7714 2070
rect 694 626 1746 628
rect 2668 626 2744 2026
rect 2988 1900 4694 2026
rect 2988 1866 3002 1900
rect 4676 1866 4694 1900
rect 2988 1852 4694 1866
rect 5768 2010 6152 2030
rect 6210 2028 7714 2036
rect 6210 2026 6722 2028
rect 6220 2022 6722 2026
rect 7500 2024 7714 2028
rect 3086 1786 4588 1852
rect 2982 1724 3054 1758
rect 3086 1752 3101 1786
rect 4577 1752 4588 1786
rect 3086 1736 4588 1752
rect 4630 1736 4934 1756
rect 2982 756 3008 1724
rect 3042 756 3054 1724
rect 2982 740 3054 756
rect 4630 1724 5054 1736
rect 4630 756 4636 1724
rect 4670 1702 5054 1724
rect 5768 1702 6110 2010
rect 4670 1042 6110 1702
rect 6144 1042 6152 2010
rect 4670 1010 6152 1042
rect 6218 1020 6340 1024
rect 7472 1020 7712 1024
rect 6210 1012 7712 1020
rect 4670 756 4994 1010
rect 6210 978 6221 1012
rect 7697 978 7712 1012
rect 6210 970 7712 978
rect 4630 746 4994 756
rect 4584 740 4994 746
rect 2982 732 4994 740
rect 5558 736 5962 738
rect 6204 736 7712 970
rect 2982 728 4680 732
rect 2982 694 3101 728
rect 4577 694 4680 728
rect 2982 682 4680 694
rect 2982 658 4604 682
rect 694 602 2784 626
rect 694 600 2244 602
rect 694 598 1268 600
rect 694 560 794 598
rect 840 594 1036 598
rect 840 560 916 594
rect 694 556 916 560
rect 962 560 1036 594
rect 1082 594 1268 598
rect 1082 560 1158 594
rect 962 556 1158 560
rect 1204 562 1268 594
rect 1314 598 2116 600
rect 1314 596 1750 598
rect 1314 562 1378 596
rect 1204 558 1378 562
rect 1424 558 1500 596
rect 1546 558 1632 596
rect 1678 560 1750 596
rect 1798 560 1874 598
rect 1922 560 2000 598
rect 2048 562 2116 598
rect 2164 564 2244 600
rect 2292 600 2784 602
rect 2292 596 2514 600
rect 2292 564 2376 596
rect 2164 562 2376 564
rect 2048 560 2376 562
rect 1678 558 2376 560
rect 2424 562 2514 596
rect 2562 596 2784 600
rect 2562 562 2616 596
rect 2424 558 2616 562
rect 2664 558 2784 596
rect 1204 556 2784 558
rect 694 526 2784 556
rect 694 524 776 526
rect 694 520 764 524
rect 1118 378 1518 526
rect 1728 524 2784 526
rect 1118 344 1132 378
rect 1506 344 1518 378
rect 1118 332 1518 344
rect 2092 370 2488 524
rect 2092 336 2102 370
rect 2476 336 2488 370
rect 1220 264 1420 332
rect 2092 322 2488 336
rect 886 220 1180 236
rect 886 186 1138 220
rect 1172 186 1180 220
rect 1220 230 1231 264
rect 1407 230 1420 264
rect 2188 256 2390 322
rect 1220 216 1420 230
rect 1812 212 2158 230
rect 2188 222 2201 256
rect 2377 222 2390 256
rect 2188 214 2390 222
rect 2720 226 2784 524
rect 3484 250 3576 658
rect 5558 546 8418 736
rect 5558 518 5962 546
rect 5558 484 5568 518
rect 5942 484 5962 518
rect 5558 466 5962 484
rect 8004 532 8418 546
rect 9060 618 9144 2308
rect 9396 2206 11592 2310
rect 11856 2298 14386 2310
rect 9396 2172 9402 2206
rect 11576 2172 11592 2206
rect 9396 2158 11592 2172
rect 11962 2204 14172 2298
rect 11962 2170 11976 2204
rect 14150 2170 14172 2204
rect 9488 2092 11494 2158
rect 11962 2146 14172 2170
rect 9488 2058 9501 2092
rect 11477 2058 11494 2092
rect 9488 2046 11494 2058
rect 12056 2090 14062 2146
rect 12056 2056 12075 2090
rect 14051 2056 14062 2090
rect 12056 2048 14062 2056
rect 9376 2044 9418 2046
rect 9344 2040 9430 2044
rect 9228 2032 9430 2040
rect 12056 2038 14056 2048
rect 9228 1880 9384 2032
rect 9228 1738 9274 1880
rect 9356 1738 9384 1880
rect 9228 1664 9384 1738
rect 9418 1664 9430 2032
rect 14096 2028 14206 2052
rect 14096 1700 14110 2028
rect 9228 1642 9430 1664
rect 14018 1660 14110 1700
rect 14144 1660 14206 2028
rect 14018 1646 14206 1660
rect 9486 1634 11492 1646
rect 9486 1600 9501 1634
rect 11477 1600 11492 1634
rect 9486 1294 11492 1600
rect 12060 1632 14206 1646
rect 12060 1598 12075 1632
rect 14051 1598 14206 1632
rect 12060 1536 14206 1598
rect 12060 1522 14172 1536
rect 12060 1294 14068 1522
rect 9486 1150 14120 1294
rect 9486 1002 10104 1150
rect 10268 1002 14120 1150
rect 9486 968 14120 1002
rect 9492 966 14120 968
rect 11164 908 14120 966
rect 11166 838 14120 908
rect 11166 672 13154 838
rect 11166 638 11172 672
rect 13148 638 13154 672
rect 11166 626 13154 638
rect 11170 624 13154 626
rect 10674 618 11102 620
rect 9060 604 11102 618
rect 9060 570 11062 604
rect 11096 570 11102 604
rect 9060 546 11102 570
rect 11166 566 13160 568
rect 11160 558 13166 566
rect 9060 542 10926 546
rect 8004 498 8020 532
rect 8394 498 8418 532
rect 8004 482 8418 498
rect 11160 524 11174 558
rect 13150 524 13166 558
rect 5652 404 5856 466
rect 5652 370 5667 404
rect 5843 370 5856 404
rect 5652 354 5856 370
rect 6072 384 6498 430
rect 6072 356 6194 384
rect 5894 342 6194 356
rect 5894 304 5902 342
rect 5936 304 6194 342
rect 886 170 1180 186
rect 1222 176 1414 188
rect 886 -46 972 170
rect 1222 142 1231 176
rect 1407 142 1414 176
rect 886 -144 974 -46
rect 558 -150 974 -144
rect 292 -218 974 -150
rect 1222 -130 1414 142
rect 1812 178 2108 212
rect 2142 178 2158 212
rect 2720 206 3454 226
rect 3484 216 3498 250
rect 3558 216 3576 250
rect 3484 206 3576 216
rect 5654 276 5858 292
rect 5894 284 6194 304
rect 5654 242 5667 276
rect 5843 242 5858 276
rect 6072 276 6194 284
rect 6306 276 6498 384
rect 8104 418 8310 482
rect 11160 458 13166 524
rect 11080 456 13250 458
rect 8104 384 8119 418
rect 8295 384 8310 418
rect 11078 444 13250 456
rect 11078 410 11084 444
rect 13240 410 13250 444
rect 8104 380 8310 384
rect 8112 374 8304 380
rect 8544 378 10392 396
rect 8544 376 10168 378
rect 8388 372 10168 376
rect 8346 356 10168 372
rect 8346 318 8354 356
rect 8388 318 10168 356
rect 8346 300 10168 318
rect 10262 300 10392 378
rect 11078 374 13250 410
rect 6072 246 6498 276
rect 8106 290 8310 300
rect 8544 290 10392 300
rect 8106 256 8119 290
rect 8295 256 8310 290
rect 1812 154 2158 178
rect 2188 168 2392 182
rect 1812 -130 1882 154
rect 1222 -162 1882 -130
rect 2188 134 2201 168
rect 2377 134 2392 168
rect 2720 172 3414 206
rect 3448 172 3454 206
rect 2720 156 3454 172
rect 3482 162 3572 174
rect 2188 -140 2392 134
rect 3482 128 3498 162
rect 3558 128 3572 162
rect 3482 64 3572 128
rect 5654 126 5858 242
rect 5652 94 5858 126
rect 3392 48 3660 64
rect 3392 14 3408 48
rect 3648 14 3660 48
rect 292 -448 382 -218
rect -26 -476 258 -472
rect -26 -536 -8 -476
rect 54 -492 258 -476
rect 292 -482 306 -448
rect 366 -482 382 -448
rect 292 -490 382 -482
rect 886 -464 974 -218
rect 1268 -204 1882 -162
rect 1268 -440 1400 -204
rect 886 -484 1238 -464
rect 1268 -474 1282 -440
rect 1388 -474 1400 -440
rect 1268 -480 1400 -474
rect 1812 -466 1882 -204
rect 2250 -202 2384 -140
rect 3392 -160 3660 14
rect 5652 -150 5856 94
rect 5652 -152 6916 -150
rect 4698 -154 6916 -152
rect 3920 -160 4000 -158
rect 3136 -170 4008 -160
rect 2250 -276 2752 -202
rect 3132 -250 4008 -170
rect 2250 -436 2384 -276
rect 1812 -480 2220 -466
rect 54 -526 208 -492
rect 242 -526 258 -492
rect 886 -518 1198 -484
rect 1232 -518 1238 -484
rect 1812 -514 2178 -480
rect 2212 -514 2220 -480
rect 2250 -470 2262 -436
rect 2368 -470 2384 -436
rect 2250 -482 2384 -470
rect 2652 -456 2750 -276
rect 3132 -430 3218 -250
rect 3920 -422 4008 -250
rect 2652 -474 3096 -456
rect 3132 -464 3142 -430
rect 3202 -464 3218 -430
rect 3132 -472 3218 -464
rect 2652 -508 3044 -474
rect 3078 -508 3096 -474
rect 3138 -476 3218 -472
rect 3442 -450 3518 -422
rect 3442 -452 3886 -450
rect 54 -536 258 -526
rect -26 -546 258 -536
rect 288 -536 382 -524
rect 886 -534 1238 -518
rect 1268 -528 1402 -516
rect 1812 -528 2220 -514
rect 2250 -514 2380 -510
rect 2250 -524 2382 -514
rect 288 -570 306 -536
rect 366 -570 382 -536
rect 288 -636 382 -570
rect 1268 -562 1282 -528
rect 1388 -562 1402 -528
rect 1268 -632 1402 -562
rect 2250 -558 2262 -524
rect 2368 -558 2382 -524
rect 2652 -524 3096 -508
rect 3126 -518 3216 -506
rect 3442 -508 3454 -452
rect 3508 -464 3886 -452
rect 3508 -498 3838 -464
rect 3872 -498 3886 -464
rect 3920 -456 3932 -422
rect 3992 -456 4008 -422
rect 3920 -466 4008 -456
rect 4698 -238 5178 -154
rect 5268 -158 6916 -154
rect 5268 -238 6294 -158
rect 4698 -242 6294 -238
rect 6384 -242 6916 -158
rect 4698 -398 6916 -242
rect 4698 -414 5700 -398
rect 4698 -448 4710 -414
rect 5686 -448 5700 -414
rect 4698 -458 5700 -448
rect 5914 -414 6916 -398
rect 8106 -372 8310 256
rect 11080 150 13250 374
rect 11020 -108 13422 150
rect 11020 -142 11030 -108
rect 13406 -142 13422 -108
rect 11020 -148 13422 -142
rect 10820 -154 10992 -152
rect 10598 -170 10992 -154
rect 11020 -158 13396 -148
rect 10598 -326 10946 -170
rect 8106 -400 8346 -372
rect 9030 -400 10042 -388
rect 5914 -448 5928 -414
rect 6904 -448 6916 -414
rect 5914 -456 6916 -448
rect 7724 -412 10042 -400
rect 7724 -446 7828 -412
rect 8804 -446 9046 -412
rect 10022 -446 10042 -412
rect 7724 -458 10042 -446
rect 6946 -462 10042 -458
rect 10598 -462 10646 -326
rect 10776 -462 10946 -326
rect 5732 -476 5886 -462
rect 3508 -508 3886 -498
rect 3924 -502 4004 -498
rect 3442 -516 3886 -508
rect 3920 -510 4004 -502
rect 2652 -526 2750 -524
rect 2250 -626 2382 -558
rect 3126 -552 3142 -518
rect 3202 -552 3216 -518
rect 3126 -614 3216 -552
rect 3920 -544 3932 -510
rect 3992 -544 4004 -510
rect 3920 -608 4004 -544
rect 5732 -544 5742 -476
rect 5776 -544 5838 -476
rect 5872 -544 5886 -476
rect 5732 -556 5886 -544
rect 6946 -474 7786 -462
rect 6946 -476 7744 -474
rect 6946 -544 6954 -476
rect 6988 -542 7744 -476
rect 7778 -542 7786 -474
rect 6988 -544 7786 -542
rect 4698 -572 5698 -562
rect 4698 -606 4710 -572
rect 5686 -606 5698 -572
rect 200 -650 466 -636
rect 200 -684 216 -650
rect 456 -684 466 -650
rect -186 -840 -150 -838
rect 200 -840 466 -684
rect 1172 -642 1490 -632
rect 1172 -676 1192 -642
rect 1478 -676 1490 -642
rect 1172 -836 1490 -676
rect 2154 -638 2470 -626
rect 2154 -672 2172 -638
rect 2458 -672 2470 -638
rect 2154 -834 2470 -672
rect 3038 -632 3308 -614
rect 3038 -666 3052 -632
rect 3292 -666 3308 -632
rect 1790 -836 2648 -834
rect 3038 -836 3308 -666
rect 3832 -624 4096 -608
rect 3832 -658 3842 -624
rect 4082 -658 4096 -624
rect 3832 -836 4096 -658
rect 4698 -668 5698 -606
rect 5918 -572 6918 -558
rect 6946 -562 7786 -544
rect 8844 -474 9006 -462
rect 8844 -542 8854 -474
rect 8888 -542 8962 -474
rect 8996 -542 9006 -474
rect 8844 -556 9006 -542
rect 10598 -538 10946 -462
rect 10980 -538 10992 -170
rect 10598 -554 10992 -538
rect 11022 -560 13412 -550
rect 5918 -606 5928 -572
rect 6904 -606 6918 -572
rect 4606 -676 5760 -668
rect 5918 -676 6918 -606
rect 7816 -570 8816 -560
rect 7816 -604 7828 -570
rect 8804 -604 8816 -570
rect 7816 -674 8816 -604
rect 9034 -570 10034 -560
rect 9034 -604 9046 -570
rect 10022 -604 10034 -570
rect 9034 -674 10034 -604
rect 11020 -566 13420 -560
rect 11020 -600 11030 -566
rect 13406 -600 13420 -566
rect 11020 -660 13420 -600
rect 7726 -676 10118 -674
rect 4606 -686 7010 -676
rect 4606 -720 4620 -686
rect 6994 -720 7010 -686
rect 4606 -834 7010 -720
rect 7726 -684 10126 -676
rect 7726 -718 7738 -684
rect 10112 -718 10126 -684
rect 7726 -832 10126 -718
rect 10934 -680 13510 -660
rect 10934 -714 10940 -680
rect 13496 -714 13510 -680
rect 10934 -824 13510 -714
rect 10626 -832 13652 -824
rect 7726 -834 13652 -832
rect 4606 -836 13652 -834
rect 766 -840 13652 -836
rect -186 -856 13652 -840
rect -186 -862 11586 -856
rect -186 -866 10790 -862
rect -186 -870 10606 -866
rect -186 -874 4638 -870
rect -186 -880 2690 -874
rect -186 -882 178 -880
rect -186 -928 -130 -882
rect -82 -928 20 -882
rect 68 -926 178 -882
rect 226 -882 710 -880
rect 226 -926 326 -882
rect 68 -928 326 -926
rect 374 -928 476 -882
rect 524 -928 622 -882
rect 670 -928 710 -882
rect 756 -884 976 -880
rect 756 -928 838 -884
rect -186 -932 838 -928
rect 888 -928 976 -884
rect 1026 -882 1548 -880
rect 1026 -928 1118 -882
rect 888 -930 1118 -928
rect 1168 -886 1406 -882
rect 1168 -930 1260 -886
rect 888 -932 1260 -930
rect -186 -934 1260 -932
rect 1310 -930 1406 -886
rect 1456 -928 1548 -882
rect 1598 -928 1720 -880
rect 1770 -882 2690 -880
rect 1770 -884 2040 -882
rect 1770 -928 1886 -884
rect 1456 -930 1886 -928
rect 1310 -932 1886 -930
rect 1940 -930 2040 -884
rect 2094 -930 2188 -882
rect 2242 -930 2330 -882
rect 2384 -930 2500 -882
rect 2554 -928 2690 -882
rect 2748 -928 2858 -874
rect 2916 -928 3030 -874
rect 3088 -928 3208 -874
rect 3266 -876 4060 -874
rect 3266 -928 3380 -876
rect 2554 -930 3380 -928
rect 3438 -880 3730 -876
rect 3438 -930 3546 -880
rect 1940 -932 3546 -930
rect 1310 -934 3546 -932
rect 3604 -930 3730 -880
rect 3788 -930 3900 -876
rect 3958 -928 4060 -876
rect 4118 -928 4240 -874
rect 4298 -876 4638 -874
rect 4298 -924 4384 -876
rect 4436 -924 4508 -876
rect 4560 -918 4638 -876
rect 4690 -918 4776 -870
rect 4828 -918 4912 -870
rect 4964 -918 5054 -870
rect 5106 -876 5542 -870
rect 5106 -918 5212 -876
rect 4560 -924 5212 -918
rect 5264 -924 5380 -876
rect 5432 -918 5542 -876
rect 5594 -872 5992 -870
rect 5594 -876 5836 -872
rect 5594 -918 5682 -876
rect 5432 -924 5682 -918
rect 5734 -920 5836 -876
rect 5888 -918 5992 -872
rect 6044 -872 10606 -870
rect 6044 -876 6284 -872
rect 6044 -918 6142 -876
rect 5888 -920 6142 -918
rect 5734 -924 6142 -920
rect 6194 -920 6284 -876
rect 6336 -920 6432 -872
rect 6484 -876 10454 -872
rect 6484 -920 6576 -876
rect 6194 -924 6576 -920
rect 6628 -924 6710 -876
rect 6762 -878 7532 -876
rect 6762 -882 7230 -878
rect 6762 -924 6840 -882
rect 4298 -928 6840 -924
rect 3958 -930 6840 -928
rect 6892 -930 6958 -882
rect 7010 -930 7092 -882
rect 7144 -926 7230 -882
rect 7282 -926 7376 -878
rect 7428 -924 7532 -878
rect 7584 -924 7702 -876
rect 7754 -880 7998 -876
rect 7754 -924 7860 -880
rect 7428 -926 7860 -924
rect 7144 -928 7860 -926
rect 7912 -924 7998 -880
rect 8050 -878 9264 -876
rect 8050 -924 8142 -878
rect 7912 -926 8142 -924
rect 8194 -880 9264 -878
rect 8194 -926 8298 -880
rect 7912 -928 8298 -926
rect 8350 -928 8434 -880
rect 8486 -928 8576 -880
rect 8628 -886 8928 -880
rect 8628 -928 8724 -886
rect 7144 -930 8724 -928
rect 3604 -934 8724 -930
rect 8776 -928 8928 -886
rect 8980 -886 9264 -880
rect 8980 -928 9100 -886
rect 8776 -934 9100 -928
rect 9152 -924 9264 -886
rect 9316 -924 9462 -876
rect 9514 -878 9934 -876
rect 9514 -880 9768 -878
rect 9514 -924 9630 -880
rect 9152 -928 9630 -924
rect 9682 -926 9768 -880
rect 9820 -924 9934 -878
rect 9986 -878 10454 -876
rect 9986 -924 10128 -878
rect 9820 -926 10128 -924
rect 10180 -882 10454 -878
rect 10180 -926 10290 -882
rect 9682 -928 10290 -926
rect 9152 -930 10290 -928
rect 10342 -930 10454 -882
rect 9152 -934 10454 -930
rect -186 -936 10454 -934
rect 10514 -930 10606 -872
rect 10666 -926 10790 -866
rect 10850 -926 11000 -862
rect 11060 -926 11196 -862
rect 11256 -926 11386 -862
rect 11446 -920 11586 -862
rect 11646 -862 13652 -856
rect 11646 -866 11946 -862
rect 11646 -920 11770 -866
rect 11446 -926 11770 -920
rect 10666 -930 11770 -926
rect 11830 -926 11946 -866
rect 12006 -866 12950 -862
rect 12006 -872 12330 -866
rect 12006 -926 12116 -872
rect 11830 -930 12116 -926
rect 10514 -936 12116 -930
rect 12176 -930 12330 -872
rect 12390 -930 12526 -866
rect 12586 -876 12950 -866
rect 12586 -930 12710 -876
rect 12176 -936 12710 -930
rect -186 -940 12710 -936
rect 12770 -926 12950 -876
rect 13010 -866 13432 -862
rect 13010 -926 13174 -866
rect 12770 -930 13174 -926
rect 13234 -926 13432 -866
rect 13492 -926 13652 -862
rect 13234 -930 13652 -926
rect 12770 -940 13652 -930
rect -186 -974 13652 -940
rect 2598 -976 13652 -974
rect 2598 -978 9278 -976
rect 2598 -980 6084 -978
rect 10626 -984 13652 -976
<< via1 >>
rect 9274 1738 9356 1880
rect 10104 1002 10268 1150
rect 6194 276 6306 384
rect 10168 300 10262 378
rect -8 -536 54 -476
rect 3454 -508 3508 -452
rect 5178 -238 5268 -154
rect 6294 -242 6384 -158
rect 10646 -462 10776 -326
<< metal2 >>
rect 6364 1880 9400 2038
rect 6364 1738 9274 1880
rect 9356 1738 9400 1880
rect 6364 1632 9400 1738
rect 6368 430 6656 1632
rect 10076 1150 10330 1190
rect 10076 1002 10104 1150
rect 10268 1002 10330 1150
rect 10076 978 10330 1002
rect 10076 842 10332 978
rect 6072 384 6656 430
rect 6072 276 6194 384
rect 6306 276 6656 384
rect 6072 246 6656 276
rect 10084 378 10332 842
rect 10084 300 10168 378
rect 10262 300 10332 378
rect 10084 250 10332 300
rect 6368 242 6656 246
rect 2060 -154 3522 -152
rect 6890 -154 10750 -152
rect -12 -238 5178 -154
rect 5268 -158 10790 -154
rect 5268 -238 6294 -158
rect -12 -242 6294 -238
rect 6384 -242 10790 -158
rect -12 -244 3522 -242
rect -12 -476 72 -244
rect -12 -536 -8 -476
rect 54 -536 72 -476
rect 3436 -452 3522 -244
rect 6890 -244 10790 -242
rect 6890 -246 10110 -244
rect 3436 -508 3454 -452
rect 3508 -508 3522 -452
rect 10636 -326 10790 -244
rect 10636 -462 10646 -326
rect 10776 -462 10790 -326
rect 10636 -476 10790 -462
rect 3436 -518 3522 -508
rect -12 -542 72 -536
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_0
timestamp 1606502482
transform 0 1 1319 -1 0 203
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_lvt_WWB6XF  sky130_fd_pr__nfet_01v8_lvt_WWB6XF_0
timestamp 1606502482
transform 0 1 336 -1 0 -509
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_RKFZUM  sky130_fd_pr__nfet_01v8_RKFZUM_0
timestamp 1606505005
transform 0 1 1335 -1 0 -501
box -211 -275 211 275
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_1
timestamp 1606502482
transform 0 1 2289 -1 0 195
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_RKFZUM  sky130_fd_pr__nfet_01v8_RKFZUM_1
timestamp 1606505005
transform 0 1 2315 -1 0 -497
box -211 -275 211 275
use sky130_fd_pr__pfet_01v8_lvt_XZ6TRL  sky130_fd_pr__pfet_01v8_lvt_XZ6TRL_0
timestamp 1606545195
transform 0 1 3839 -1 0 1240
box -696 -969 696 969
use sky130_fd_pr__nfet_01v8_WWB6XF  sky130_fd_pr__nfet_01v8_WWB6XF_0
timestamp 1606508276
transform 0 1 3172 -1 0 -491
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_WWB6XF  sky130_fd_pr__nfet_01v8_WWB6XF_1
timestamp 1606508276
transform 0 1 3962 -1 0 -483
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_WWB6XF  sky130_fd_pr__nfet_01v8_WWB6XF_2
timestamp 1606508276
transform 0 1 3528 -1 0 189
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_XAABVK  sky130_fd_pr__nfet_01v8_XAABVK_0
timestamp 1606545195
transform 0 1 5807 -1 0 -510
box -246 -1319 246 1319
use sky130_fd_pr__pfet_01v8_lvt_2CKJF2  sky130_fd_pr__pfet_01v8_lvt_2CKJF2_0
timestamp 1606545195
transform 0 1 5755 -1 0 323
box -231 -319 231 319
use sky130_fd_pr__pfet_01v8_lvt_2CKJF2  sky130_fd_pr__pfet_01v8_lvt_2CKJF2_1
timestamp 1606545195
transform 0 1 8207 -1 0 337
box -231 -319 231 319
use sky130_fd_pr__nfet_01v8_XAABVK  sky130_fd_pr__nfet_01v8_XAABVK_1
timestamp 1606545195
transform 0 1 8925 -1 0 -508
box -246 -1319 246 1319
use sky130_fd_pr__nfet_01v8_lvt_6NXDEK  sky130_fd_pr__nfet_01v8_lvt_6NXDEK_0
timestamp 1606601234
transform 0 1 12162 -1 0 585
box -211 -1210 211 1210
use sky130_fd_pr__nfet_01v8_lvt_VCXMU2  sky130_fd_pr__nfet_01v8_lvt_VCXMU2_0
timestamp 1606601234
transform 0 1 12218 -1 0 -354
box -396 -1410 396 1410
use sky130_fd_pr__pfet_01v8_lvt_XZ6TRL  sky130_fd_pr__pfet_01v8_lvt_XZ6TRL_1
timestamp 1606545195
transform 0 1 6959 -1 0 1524
box -696 -969 696 969
use sky130_fd_pr__pfet_01v8_lvt_ZJ2V3W  sky130_fd_pr__pfet_01v8_lvt_ZJ2V3W_1
timestamp 1606606258
transform 0 1 13063 -1 0 1844
box -396 -1219 396 1219
use sky130_fd_pr__pfet_01v8_lvt_ZJ2V3W  sky130_fd_pr__pfet_01v8_lvt_ZJ2V3W_0
timestamp 1606606258
transform 0 1 10489 -1 0 1846
box -396 -1219 396 1219
<< labels >>
rlabel metal1 302 -224 366 -156 1 Inv1IN
port 2 n
rlabel metal1 304 -932 368 -864 1 Gnd
port 4 n
rlabel metal1 1284 -204 1372 -146 1 Inv2IN
port 5 n
rlabel metal1 2272 -214 2370 -116 1 Vinit
port 6 n
rlabel metal1 3504 -124 3562 -60 1 AmpBias2
port 7 n
rlabel metal1 6084 296 6130 348 1 Vcntrl
port 8 n
rlabel metal1 8576 304 8634 364 1 DiifAmpPos
port 9 n
rlabel via1 0 -530 48 -486 1 vbn
port 1 n
<< end >>
