magic
tech sky130A
magscale 1 2
timestamp 1606057846
<< nwell >>
rect -1352 -1219 1352 1219
<< pmos >>
rect -1156 -1000 -1056 1000
rect -998 -1000 -898 1000
rect -840 -1000 -740 1000
rect -682 -1000 -582 1000
rect -524 -1000 -424 1000
rect -366 -1000 -266 1000
rect -208 -1000 -108 1000
rect -50 -1000 50 1000
rect 108 -1000 208 1000
rect 266 -1000 366 1000
rect 424 -1000 524 1000
rect 582 -1000 682 1000
rect 740 -1000 840 1000
rect 898 -1000 998 1000
rect 1056 -1000 1156 1000
<< pdiff >>
rect -1214 988 -1156 1000
rect -1214 -988 -1202 988
rect -1168 -988 -1156 988
rect -1214 -1000 -1156 -988
rect -1056 988 -998 1000
rect -1056 -988 -1044 988
rect -1010 -988 -998 988
rect -1056 -1000 -998 -988
rect -898 988 -840 1000
rect -898 -988 -886 988
rect -852 -988 -840 988
rect -898 -1000 -840 -988
rect -740 988 -682 1000
rect -740 -988 -728 988
rect -694 -988 -682 988
rect -740 -1000 -682 -988
rect -582 988 -524 1000
rect -582 -988 -570 988
rect -536 -988 -524 988
rect -582 -1000 -524 -988
rect -424 988 -366 1000
rect -424 -988 -412 988
rect -378 -988 -366 988
rect -424 -1000 -366 -988
rect -266 988 -208 1000
rect -266 -988 -254 988
rect -220 -988 -208 988
rect -266 -1000 -208 -988
rect -108 988 -50 1000
rect -108 -988 -96 988
rect -62 -988 -50 988
rect -108 -1000 -50 -988
rect 50 988 108 1000
rect 50 -988 62 988
rect 96 -988 108 988
rect 50 -1000 108 -988
rect 208 988 266 1000
rect 208 -988 220 988
rect 254 -988 266 988
rect 208 -1000 266 -988
rect 366 988 424 1000
rect 366 -988 378 988
rect 412 -988 424 988
rect 366 -1000 424 -988
rect 524 988 582 1000
rect 524 -988 536 988
rect 570 -988 582 988
rect 524 -1000 582 -988
rect 682 988 740 1000
rect 682 -988 694 988
rect 728 -988 740 988
rect 682 -1000 740 -988
rect 840 988 898 1000
rect 840 -988 852 988
rect 886 -988 898 988
rect 840 -1000 898 -988
rect 998 988 1056 1000
rect 998 -988 1010 988
rect 1044 -988 1056 988
rect 998 -1000 1056 -988
rect 1156 988 1214 1000
rect 1156 -988 1168 988
rect 1202 -988 1214 988
rect 1156 -1000 1214 -988
<< pdiffc >>
rect -1202 -988 -1168 988
rect -1044 -988 -1010 988
rect -886 -988 -852 988
rect -728 -988 -694 988
rect -570 -988 -536 988
rect -412 -988 -378 988
rect -254 -988 -220 988
rect -96 -988 -62 988
rect 62 -988 96 988
rect 220 -988 254 988
rect 378 -988 412 988
rect 536 -988 570 988
rect 694 -988 728 988
rect 852 -988 886 988
rect 1010 -988 1044 988
rect 1168 -988 1202 988
<< nsubdiff >>
rect -1316 1149 -1220 1183
rect 1220 1149 1316 1183
rect -1316 1087 -1282 1149
rect 1282 1087 1316 1149
rect -1316 -1149 -1282 -1087
rect 1282 -1149 1316 -1087
rect -1316 -1183 -1220 -1149
rect 1220 -1183 1316 -1149
<< nsubdiffcont >>
rect -1220 1149 1220 1183
rect -1316 -1087 -1282 1087
rect 1282 -1087 1316 1087
rect -1220 -1183 1220 -1149
<< poly >>
rect -1156 1081 -1056 1097
rect -1156 1047 -1140 1081
rect -1072 1047 -1056 1081
rect -1156 1000 -1056 1047
rect -998 1081 -898 1097
rect -998 1047 -982 1081
rect -914 1047 -898 1081
rect -998 1000 -898 1047
rect -840 1081 -740 1097
rect -840 1047 -824 1081
rect -756 1047 -740 1081
rect -840 1000 -740 1047
rect -682 1081 -582 1097
rect -682 1047 -666 1081
rect -598 1047 -582 1081
rect -682 1000 -582 1047
rect -524 1081 -424 1097
rect -524 1047 -508 1081
rect -440 1047 -424 1081
rect -524 1000 -424 1047
rect -366 1081 -266 1097
rect -366 1047 -350 1081
rect -282 1047 -266 1081
rect -366 1000 -266 1047
rect -208 1081 -108 1097
rect -208 1047 -192 1081
rect -124 1047 -108 1081
rect -208 1000 -108 1047
rect -50 1081 50 1097
rect -50 1047 -34 1081
rect 34 1047 50 1081
rect -50 1000 50 1047
rect 108 1081 208 1097
rect 108 1047 124 1081
rect 192 1047 208 1081
rect 108 1000 208 1047
rect 266 1081 366 1097
rect 266 1047 282 1081
rect 350 1047 366 1081
rect 266 1000 366 1047
rect 424 1081 524 1097
rect 424 1047 440 1081
rect 508 1047 524 1081
rect 424 1000 524 1047
rect 582 1081 682 1097
rect 582 1047 598 1081
rect 666 1047 682 1081
rect 582 1000 682 1047
rect 740 1081 840 1097
rect 740 1047 756 1081
rect 824 1047 840 1081
rect 740 1000 840 1047
rect 898 1081 998 1097
rect 898 1047 914 1081
rect 982 1047 998 1081
rect 898 1000 998 1047
rect 1056 1081 1156 1097
rect 1056 1047 1072 1081
rect 1140 1047 1156 1081
rect 1056 1000 1156 1047
rect -1156 -1047 -1056 -1000
rect -1156 -1081 -1140 -1047
rect -1072 -1081 -1056 -1047
rect -1156 -1097 -1056 -1081
rect -998 -1047 -898 -1000
rect -998 -1081 -982 -1047
rect -914 -1081 -898 -1047
rect -998 -1097 -898 -1081
rect -840 -1047 -740 -1000
rect -840 -1081 -824 -1047
rect -756 -1081 -740 -1047
rect -840 -1097 -740 -1081
rect -682 -1047 -582 -1000
rect -682 -1081 -666 -1047
rect -598 -1081 -582 -1047
rect -682 -1097 -582 -1081
rect -524 -1047 -424 -1000
rect -524 -1081 -508 -1047
rect -440 -1081 -424 -1047
rect -524 -1097 -424 -1081
rect -366 -1047 -266 -1000
rect -366 -1081 -350 -1047
rect -282 -1081 -266 -1047
rect -366 -1097 -266 -1081
rect -208 -1047 -108 -1000
rect -208 -1081 -192 -1047
rect -124 -1081 -108 -1047
rect -208 -1097 -108 -1081
rect -50 -1047 50 -1000
rect -50 -1081 -34 -1047
rect 34 -1081 50 -1047
rect -50 -1097 50 -1081
rect 108 -1047 208 -1000
rect 108 -1081 124 -1047
rect 192 -1081 208 -1047
rect 108 -1097 208 -1081
rect 266 -1047 366 -1000
rect 266 -1081 282 -1047
rect 350 -1081 366 -1047
rect 266 -1097 366 -1081
rect 424 -1047 524 -1000
rect 424 -1081 440 -1047
rect 508 -1081 524 -1047
rect 424 -1097 524 -1081
rect 582 -1047 682 -1000
rect 582 -1081 598 -1047
rect 666 -1081 682 -1047
rect 582 -1097 682 -1081
rect 740 -1047 840 -1000
rect 740 -1081 756 -1047
rect 824 -1081 840 -1047
rect 740 -1097 840 -1081
rect 898 -1047 998 -1000
rect 898 -1081 914 -1047
rect 982 -1081 998 -1047
rect 898 -1097 998 -1081
rect 1056 -1047 1156 -1000
rect 1056 -1081 1072 -1047
rect 1140 -1081 1156 -1047
rect 1056 -1097 1156 -1081
<< polycont >>
rect -1140 1047 -1072 1081
rect -982 1047 -914 1081
rect -824 1047 -756 1081
rect -666 1047 -598 1081
rect -508 1047 -440 1081
rect -350 1047 -282 1081
rect -192 1047 -124 1081
rect -34 1047 34 1081
rect 124 1047 192 1081
rect 282 1047 350 1081
rect 440 1047 508 1081
rect 598 1047 666 1081
rect 756 1047 824 1081
rect 914 1047 982 1081
rect 1072 1047 1140 1081
rect -1140 -1081 -1072 -1047
rect -982 -1081 -914 -1047
rect -824 -1081 -756 -1047
rect -666 -1081 -598 -1047
rect -508 -1081 -440 -1047
rect -350 -1081 -282 -1047
rect -192 -1081 -124 -1047
rect -34 -1081 34 -1047
rect 124 -1081 192 -1047
rect 282 -1081 350 -1047
rect 440 -1081 508 -1047
rect 598 -1081 666 -1047
rect 756 -1081 824 -1047
rect 914 -1081 982 -1047
rect 1072 -1081 1140 -1047
<< locali >>
rect -1316 1149 -1220 1183
rect 1220 1149 1316 1183
rect -1316 1087 -1282 1149
rect 1282 1087 1316 1149
rect -1156 1047 -1140 1081
rect -1072 1047 -1056 1081
rect -998 1047 -982 1081
rect -914 1047 -898 1081
rect -840 1047 -824 1081
rect -756 1047 -740 1081
rect -682 1047 -666 1081
rect -598 1047 -582 1081
rect -524 1047 -508 1081
rect -440 1047 -424 1081
rect -366 1047 -350 1081
rect -282 1047 -266 1081
rect -208 1047 -192 1081
rect -124 1047 -108 1081
rect -50 1047 -34 1081
rect 34 1047 50 1081
rect 108 1047 124 1081
rect 192 1047 208 1081
rect 266 1047 282 1081
rect 350 1047 366 1081
rect 424 1047 440 1081
rect 508 1047 524 1081
rect 582 1047 598 1081
rect 666 1047 682 1081
rect 740 1047 756 1081
rect 824 1047 840 1081
rect 898 1047 914 1081
rect 982 1047 998 1081
rect 1056 1047 1072 1081
rect 1140 1047 1156 1081
rect -1202 988 -1168 1004
rect -1202 -1004 -1168 -988
rect -1044 988 -1010 1004
rect -1044 -1004 -1010 -988
rect -886 988 -852 1004
rect -886 -1004 -852 -988
rect -728 988 -694 1004
rect -728 -1004 -694 -988
rect -570 988 -536 1004
rect -570 -1004 -536 -988
rect -412 988 -378 1004
rect -412 -1004 -378 -988
rect -254 988 -220 1004
rect -254 -1004 -220 -988
rect -96 988 -62 1004
rect -96 -1004 -62 -988
rect 62 988 96 1004
rect 62 -1004 96 -988
rect 220 988 254 1004
rect 220 -1004 254 -988
rect 378 988 412 1004
rect 378 -1004 412 -988
rect 536 988 570 1004
rect 536 -1004 570 -988
rect 694 988 728 1004
rect 694 -1004 728 -988
rect 852 988 886 1004
rect 852 -1004 886 -988
rect 1010 988 1044 1004
rect 1010 -1004 1044 -988
rect 1168 988 1202 1004
rect 1168 -1004 1202 -988
rect -1156 -1081 -1140 -1047
rect -1072 -1081 -1056 -1047
rect -998 -1081 -982 -1047
rect -914 -1081 -898 -1047
rect -840 -1081 -824 -1047
rect -756 -1081 -740 -1047
rect -682 -1081 -666 -1047
rect -598 -1081 -582 -1047
rect -524 -1081 -508 -1047
rect -440 -1081 -424 -1047
rect -366 -1081 -350 -1047
rect -282 -1081 -266 -1047
rect -208 -1081 -192 -1047
rect -124 -1081 -108 -1047
rect -50 -1081 -34 -1047
rect 34 -1081 50 -1047
rect 108 -1081 124 -1047
rect 192 -1081 208 -1047
rect 266 -1081 282 -1047
rect 350 -1081 366 -1047
rect 424 -1081 440 -1047
rect 508 -1081 524 -1047
rect 582 -1081 598 -1047
rect 666 -1081 682 -1047
rect 740 -1081 756 -1047
rect 824 -1081 840 -1047
rect 898 -1081 914 -1047
rect 982 -1081 998 -1047
rect 1056 -1081 1072 -1047
rect 1140 -1081 1156 -1047
rect -1316 -1149 -1282 -1087
rect 1282 -1149 1316 -1087
rect -1316 -1183 -1220 -1149
rect 1220 -1183 1316 -1149
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1299 -1166 1299 1166
string parameters w 10 l 0.5 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
