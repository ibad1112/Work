magic
tech sky130A
timestamp 1606420870
<< pwell >>
rect -1343 -705 1343 705
<< nmoslvt >>
rect -1245 -600 -1045 600
rect -1016 -600 -816 600
rect -787 -600 -587 600
rect -558 -600 -358 600
rect -329 -600 -129 600
rect -100 -600 100 600
rect 129 -600 329 600
rect 358 -600 558 600
rect 587 -600 787 600
rect 816 -600 1016 600
rect 1045 -600 1245 600
<< ndiff >>
rect -1274 594 -1245 600
rect -1274 -594 -1268 594
rect -1251 -594 -1245 594
rect -1274 -600 -1245 -594
rect -1045 594 -1016 600
rect -1045 -594 -1039 594
rect -1022 -594 -1016 594
rect -1045 -600 -1016 -594
rect -816 594 -787 600
rect -816 -594 -810 594
rect -793 -594 -787 594
rect -816 -600 -787 -594
rect -587 594 -558 600
rect -587 -594 -581 594
rect -564 -594 -558 594
rect -587 -600 -558 -594
rect -358 594 -329 600
rect -358 -594 -352 594
rect -335 -594 -329 594
rect -358 -600 -329 -594
rect -129 594 -100 600
rect -129 -594 -123 594
rect -106 -594 -100 594
rect -129 -600 -100 -594
rect 100 594 129 600
rect 100 -594 106 594
rect 123 -594 129 594
rect 100 -600 129 -594
rect 329 594 358 600
rect 329 -594 335 594
rect 352 -594 358 594
rect 329 -600 358 -594
rect 558 594 587 600
rect 558 -594 564 594
rect 581 -594 587 594
rect 558 -600 587 -594
rect 787 594 816 600
rect 787 -594 793 594
rect 810 -594 816 594
rect 787 -600 816 -594
rect 1016 594 1045 600
rect 1016 -594 1022 594
rect 1039 -594 1045 594
rect 1016 -600 1045 -594
rect 1245 594 1274 600
rect 1245 -594 1251 594
rect 1268 -594 1274 594
rect 1245 -600 1274 -594
<< ndiffc >>
rect -1268 -594 -1251 594
rect -1039 -594 -1022 594
rect -810 -594 -793 594
rect -581 -594 -564 594
rect -352 -594 -335 594
rect -123 -594 -106 594
rect 106 -594 123 594
rect 335 -594 352 594
rect 564 -594 581 594
rect 793 -594 810 594
rect 1022 -594 1039 594
rect 1251 -594 1268 594
<< psubdiff >>
rect -1325 670 -1277 687
rect 1277 670 1325 687
rect -1325 639 -1308 670
rect 1308 639 1325 670
rect -1325 -670 -1308 -639
rect 1308 -670 1325 -639
rect -1325 -687 -1277 -670
rect 1277 -687 1325 -670
<< psubdiffcont >>
rect -1277 670 1277 687
rect -1325 -639 -1308 639
rect 1308 -639 1325 639
rect -1277 -687 1277 -670
<< poly >>
rect -1245 636 -1045 644
rect -1245 619 -1237 636
rect -1053 619 -1045 636
rect -1245 600 -1045 619
rect -1016 636 -816 644
rect -1016 619 -1008 636
rect -824 619 -816 636
rect -1016 600 -816 619
rect -787 636 -587 644
rect -787 619 -779 636
rect -595 619 -587 636
rect -787 600 -587 619
rect -558 636 -358 644
rect -558 619 -550 636
rect -366 619 -358 636
rect -558 600 -358 619
rect -329 636 -129 644
rect -329 619 -321 636
rect -137 619 -129 636
rect -329 600 -129 619
rect -100 636 100 644
rect -100 619 -92 636
rect 92 619 100 636
rect -100 600 100 619
rect 129 636 329 644
rect 129 619 137 636
rect 321 619 329 636
rect 129 600 329 619
rect 358 636 558 644
rect 358 619 366 636
rect 550 619 558 636
rect 358 600 558 619
rect 587 636 787 644
rect 587 619 595 636
rect 779 619 787 636
rect 587 600 787 619
rect 816 636 1016 644
rect 816 619 824 636
rect 1008 619 1016 636
rect 816 600 1016 619
rect 1045 636 1245 644
rect 1045 619 1053 636
rect 1237 619 1245 636
rect 1045 600 1245 619
rect -1245 -619 -1045 -600
rect -1245 -636 -1237 -619
rect -1053 -636 -1045 -619
rect -1245 -644 -1045 -636
rect -1016 -619 -816 -600
rect -1016 -636 -1008 -619
rect -824 -636 -816 -619
rect -1016 -644 -816 -636
rect -787 -619 -587 -600
rect -787 -636 -779 -619
rect -595 -636 -587 -619
rect -787 -644 -587 -636
rect -558 -619 -358 -600
rect -558 -636 -550 -619
rect -366 -636 -358 -619
rect -558 -644 -358 -636
rect -329 -619 -129 -600
rect -329 -636 -321 -619
rect -137 -636 -129 -619
rect -329 -644 -129 -636
rect -100 -619 100 -600
rect -100 -636 -92 -619
rect 92 -636 100 -619
rect -100 -644 100 -636
rect 129 -619 329 -600
rect 129 -636 137 -619
rect 321 -636 329 -619
rect 129 -644 329 -636
rect 358 -619 558 -600
rect 358 -636 366 -619
rect 550 -636 558 -619
rect 358 -644 558 -636
rect 587 -619 787 -600
rect 587 -636 595 -619
rect 779 -636 787 -619
rect 587 -644 787 -636
rect 816 -619 1016 -600
rect 816 -636 824 -619
rect 1008 -636 1016 -619
rect 816 -644 1016 -636
rect 1045 -619 1245 -600
rect 1045 -636 1053 -619
rect 1237 -636 1245 -619
rect 1045 -644 1245 -636
<< polycont >>
rect -1237 619 -1053 636
rect -1008 619 -824 636
rect -779 619 -595 636
rect -550 619 -366 636
rect -321 619 -137 636
rect -92 619 92 636
rect 137 619 321 636
rect 366 619 550 636
rect 595 619 779 636
rect 824 619 1008 636
rect 1053 619 1237 636
rect -1237 -636 -1053 -619
rect -1008 -636 -824 -619
rect -779 -636 -595 -619
rect -550 -636 -366 -619
rect -321 -636 -137 -619
rect -92 -636 92 -619
rect 137 -636 321 -619
rect 366 -636 550 -619
rect 595 -636 779 -619
rect 824 -636 1008 -619
rect 1053 -636 1237 -619
<< locali >>
rect -1325 670 -1277 687
rect 1277 670 1325 687
rect -1325 639 -1308 670
rect 1308 639 1325 670
rect -1245 619 -1237 636
rect -1053 619 -1045 636
rect -1016 619 -1008 636
rect -824 619 -816 636
rect -787 619 -779 636
rect -595 619 -587 636
rect -558 619 -550 636
rect -366 619 -358 636
rect -329 619 -321 636
rect -137 619 -129 636
rect -100 619 -92 636
rect 92 619 100 636
rect 129 619 137 636
rect 321 619 329 636
rect 358 619 366 636
rect 550 619 558 636
rect 587 619 595 636
rect 779 619 787 636
rect 816 619 824 636
rect 1008 619 1016 636
rect 1045 619 1053 636
rect 1237 619 1245 636
rect -1268 594 -1251 602
rect -1268 -602 -1251 -594
rect -1039 594 -1022 602
rect -1039 -602 -1022 -594
rect -810 594 -793 602
rect -810 -602 -793 -594
rect -581 594 -564 602
rect -581 -602 -564 -594
rect -352 594 -335 602
rect -352 -602 -335 -594
rect -123 594 -106 602
rect -123 -602 -106 -594
rect 106 594 123 602
rect 106 -602 123 -594
rect 335 594 352 602
rect 335 -602 352 -594
rect 564 594 581 602
rect 564 -602 581 -594
rect 793 594 810 602
rect 793 -602 810 -594
rect 1022 594 1039 602
rect 1022 -602 1039 -594
rect 1251 594 1268 602
rect 1251 -602 1268 -594
rect -1245 -636 -1237 -619
rect -1053 -636 -1045 -619
rect -1016 -636 -1008 -619
rect -824 -636 -816 -619
rect -787 -636 -779 -619
rect -595 -636 -587 -619
rect -558 -636 -550 -619
rect -366 -636 -358 -619
rect -329 -636 -321 -619
rect -137 -636 -129 -619
rect -100 -636 -92 -619
rect 92 -636 100 -619
rect 129 -636 137 -619
rect 321 -636 329 -619
rect 358 -636 366 -619
rect 550 -636 558 -619
rect 587 -636 595 -619
rect 779 -636 787 -619
rect 816 -636 824 -619
rect 1008 -636 1016 -619
rect 1045 -636 1053 -619
rect 1237 -636 1245 -619
rect -1325 -670 -1308 -639
rect 1308 -670 1325 -639
rect -1325 -687 -1277 -670
rect 1277 -687 1325 -670
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -1316 -678 1316 678
string parameters w 12 l 2 m 1 nf 11 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
