magic
tech sky130A
magscale 1 2
timestamp 1606606258
<< nwell >>
rect -396 -1219 396 1219
<< pmoslvt >>
rect -200 -1000 200 1000
<< pdiff >>
rect -258 988 -200 1000
rect -258 -988 -246 988
rect -212 -988 -200 988
rect -258 -1000 -200 -988
rect 200 988 258 1000
rect 200 -988 212 988
rect 246 -988 258 988
rect 200 -1000 258 -988
<< pdiffc >>
rect -246 -988 -212 988
rect 212 -988 246 988
<< nsubdiff >>
rect -360 1149 -264 1183
rect 264 1149 360 1183
rect -360 1087 -326 1149
rect 326 1087 360 1149
rect -360 -1149 -326 -1087
rect 326 -1149 360 -1087
rect -360 -1183 -264 -1149
rect 264 -1183 360 -1149
<< nsubdiffcont >>
rect -264 1149 264 1183
rect -360 -1087 -326 1087
rect 326 -1087 360 1087
rect -264 -1183 264 -1149
<< poly >>
rect -200 1081 200 1097
rect -200 1047 -184 1081
rect 184 1047 200 1081
rect -200 1000 200 1047
rect -200 -1047 200 -1000
rect -200 -1081 -184 -1047
rect 184 -1081 200 -1047
rect -200 -1097 200 -1081
<< polycont >>
rect -184 1047 184 1081
rect -184 -1081 184 -1047
<< locali >>
rect -360 1149 -264 1183
rect 264 1149 360 1183
rect -360 1087 -326 1149
rect 326 1087 360 1149
rect -200 1047 -184 1081
rect 184 1047 200 1081
rect -246 988 -212 1004
rect -246 -1004 -212 -988
rect 212 988 246 1004
rect 212 -1004 246 -988
rect -200 -1081 -184 -1047
rect 184 -1081 200 -1047
rect -360 -1149 -326 -1087
rect 326 -1149 360 -1087
rect -360 -1183 -264 -1149
rect 264 -1183 360 -1149
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -343 -1166 343 1166
string parameters w 10 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
