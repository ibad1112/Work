magic
tech sky130A
magscale 1 2
timestamp 1606420870
<< nwell >>
rect 8208 2782 10390 2790
rect 8104 2780 10390 2782
rect 7702 2774 10390 2780
rect 4886 2770 10390 2774
rect 2344 2734 10390 2770
rect -128 2350 10390 2734
rect 2042 2342 10390 2350
rect 2042 2332 3072 2342
rect 2042 -58 2844 2332
rect 4820 2326 10390 2342
rect 4820 -72 10260 2326
<< pwell >>
rect 3612 -1196 6708 -756
<< psubdiff >>
rect 3588 -4774 9120 -4720
rect 3588 -4778 7934 -4774
rect 3588 -4784 5066 -4778
rect 3588 -4900 4172 -4784
rect 4330 -4894 5066 -4784
rect 5224 -4894 6836 -4778
rect 6994 -4890 7934 -4778
rect 8092 -4890 9120 -4774
rect 6994 -4894 9120 -4890
rect 4330 -4900 9120 -4894
rect 3588 -4948 9120 -4900
<< nsubdiff >>
rect 7760 2668 10230 2688
rect 4766 2666 10230 2668
rect 2 2654 10230 2666
rect 2 2636 6052 2654
rect 2 2626 3260 2636
rect 2 2616 1418 2626
rect 2 2522 484 2616
rect 620 2532 1418 2616
rect 1554 2546 3260 2626
rect 3372 2628 6052 2636
rect 3372 2546 4178 2628
rect 1554 2538 4178 2546
rect 4290 2552 6052 2628
rect 6158 2648 10230 2654
rect 6158 2552 7014 2648
rect 4290 2546 7014 2552
rect 7120 2642 10230 2648
rect 7120 2640 9538 2642
rect 7120 2548 8592 2640
rect 8682 2550 9538 2640
rect 9628 2550 10230 2642
rect 8682 2548 10230 2550
rect 7120 2546 10230 2548
rect 4290 2538 10230 2546
rect 1554 2532 10230 2538
rect 620 2522 10230 2532
rect 2 2514 10230 2522
rect 2 2506 2124 2514
rect 4766 2510 10230 2514
rect 7760 2506 10230 2510
<< psubdiffcont >>
rect 4172 -4900 4330 -4784
rect 5066 -4894 5224 -4778
rect 6836 -4894 6994 -4778
rect 7934 -4890 8092 -4774
<< nsubdiffcont >>
rect 484 2522 620 2616
rect 1418 2532 1554 2626
rect 3260 2546 3372 2636
rect 4178 2538 4290 2628
rect 6052 2552 6158 2654
rect 7014 2546 7120 2648
rect 8592 2548 8682 2640
rect 9538 2550 9628 2642
<< locali >>
rect 8660 2662 10214 2666
rect 4726 2654 9084 2662
rect 4726 2646 6052 2654
rect 2018 2644 6052 2646
rect 2018 2642 5658 2644
rect 6 2638 5658 2642
rect 6 2636 3732 2638
rect 6 2628 3260 2636
rect 6 2626 2840 2628
rect 6 2616 1418 2626
rect 6 2604 484 2616
rect 6 2532 142 2604
rect 242 2532 484 2604
rect 6 2522 484 2532
rect 620 2612 1418 2616
rect 620 2540 978 2612
rect 1078 2540 1418 2612
rect 620 2532 1418 2540
rect 1554 2624 2840 2626
rect 1554 2552 1888 2624
rect 1988 2552 2840 2624
rect 1554 2538 2840 2552
rect 2952 2546 3260 2628
rect 3372 2548 3732 2636
rect 3844 2628 5658 2638
rect 3844 2548 4178 2628
rect 3372 2546 4178 2548
rect 2952 2538 4178 2546
rect 4290 2626 5658 2628
rect 4290 2538 4622 2626
rect 1554 2536 4622 2538
rect 4734 2542 5658 2626
rect 5764 2552 6052 2644
rect 6158 2648 8172 2654
rect 6158 2634 7014 2648
rect 6158 2552 6512 2634
rect 5764 2542 6512 2552
rect 4734 2536 6512 2542
rect 1554 2534 6512 2536
rect 1554 2532 4756 2534
rect 6618 2546 7014 2634
rect 7120 2634 8172 2648
rect 7120 2546 7472 2634
rect 6618 2534 7472 2546
rect 7578 2538 8172 2634
rect 8268 2640 9084 2654
rect 8268 2548 8592 2640
rect 8682 2548 9084 2640
rect 8268 2546 9084 2548
rect 9180 2660 10214 2662
rect 9180 2642 10012 2660
rect 9180 2550 9538 2642
rect 9628 2550 10012 2642
rect 9180 2546 10012 2550
rect 8268 2544 10012 2546
rect 10108 2544 10214 2660
rect 8268 2540 10214 2544
rect 8268 2538 8796 2540
rect 7578 2534 8796 2538
rect 620 2528 4756 2532
rect 620 2522 2116 2528
rect 8260 2206 8628 2240
rect 8718 2206 9086 2240
rect 9176 2206 9544 2240
rect 9634 2206 10002 2240
rect 3614 -4764 9092 -4762
rect 3614 -4770 6492 -4764
rect 3614 -4878 3716 -4770
rect 3830 -4778 5552 -4770
rect 3830 -4784 5066 -4778
rect 3830 -4878 4172 -4784
rect 3614 -4900 4172 -4878
rect 4330 -4786 5066 -4784
rect 4330 -4894 4662 -4786
rect 4776 -4894 5066 -4786
rect 5224 -4878 5552 -4778
rect 5666 -4872 6492 -4770
rect 6606 -4770 8314 -4764
rect 6606 -4778 7420 -4770
rect 6606 -4872 6836 -4778
rect 5666 -4878 6836 -4872
rect 5224 -4894 6836 -4878
rect 6994 -4878 7420 -4778
rect 7534 -4774 8314 -4770
rect 7534 -4878 7934 -4774
rect 6994 -4890 7934 -4878
rect 8092 -4872 8314 -4774
rect 8428 -4872 9092 -4764
rect 8092 -4890 9092 -4872
rect 6994 -4894 9092 -4890
rect 4330 -4900 9092 -4894
rect 3614 -4912 9092 -4900
<< viali >>
rect 142 2532 242 2604
rect 978 2540 1078 2612
rect 1888 2552 1988 2624
rect 2840 2538 2952 2628
rect 3732 2548 3844 2638
rect 4622 2536 4734 2626
rect 5658 2542 5764 2644
rect 6512 2532 6618 2634
rect 7472 2532 7578 2634
rect 8172 2538 8268 2654
rect 9084 2546 9180 2662
rect 10012 2544 10108 2660
rect 76 2308 148 2344
rect 3596 2322 3672 2366
rect 6100 2284 6170 2330
rect 8800 2308 8866 2352
rect 2920 2210 3288 2244
rect 3378 2210 3746 2244
rect 3836 2210 4204 2244
rect 4294 2210 4662 2244
rect 5736 2184 6104 2218
rect 6194 2184 6562 2218
rect 6652 2184 7020 2218
rect 7110 2184 7478 2218
rect 96 1978 130 2050
rect 1018 1974 1052 2046
rect 1932 1974 1966 2046
rect 2852 1980 2888 2062
rect 3770 1974 3806 2056
rect 4684 1974 4720 2056
rect 5672 1964 5722 2056
rect 6592 1966 6632 2052
rect 7504 1974 7544 2060
rect 8202 1968 8238 2030
rect 9124 1966 9162 2058
rect 10032 1976 10070 2068
rect 3310 1762 3346 1844
rect 4238 1756 4274 1838
rect 560 1664 594 1736
rect 1470 1664 1506 1742
rect 6134 1678 6174 1764
rect 7050 1678 7090 1764
rect 8636 1572 8704 1678
rect 9558 1580 9626 1686
rect 159 85 527 119
rect 617 85 985 119
rect 1075 85 1443 119
rect 1533 85 1901 119
rect 8260 78 8628 112
rect 8718 78 9086 112
rect 9176 78 9544 112
rect 9634 78 10002 112
rect 2328 -948 2468 -912
rect 7816 -940 7900 -900
rect 2362 -1054 2468 -1008
rect 7816 -1036 7896 -996
rect 2354 -1162 2460 -1116
rect 7818 -1142 7898 -1102
rect 3766 -2180 3814 -2084
rect 4682 -2188 4730 -2092
rect 5600 -2176 5648 -2080
rect 6508 -2168 6556 -2072
rect 7414 -2174 7462 -2078
rect 8346 -2174 8394 -2078
rect 4198 -2396 4268 -2286
rect 5122 -2384 5192 -2274
rect 6040 -2372 6110 -2262
rect 6964 -2372 7034 -2262
rect 7888 -2384 7958 -2274
rect 8784 -2366 8854 -2256
rect 3835 -4461 4203 -4427
rect 4293 -4461 4661 -4427
rect 4751 -4461 5119 -4427
rect 5209 -4461 5577 -4427
rect 5667 -4461 6035 -4427
rect 6125 -4461 6493 -4427
rect 6583 -4461 6951 -4427
rect 7041 -4461 7409 -4427
rect 7499 -4461 7867 -4427
rect 7957 -4461 8325 -4427
rect 8415 -4461 8783 -4427
rect 7688 -4572 7790 -4538
rect 3716 -4878 3830 -4770
rect 4662 -4894 4776 -4786
rect 5552 -4878 5666 -4770
rect 6492 -4872 6606 -4764
rect 7420 -4878 7534 -4770
rect 8314 -4872 8428 -4764
<< metal1 >>
rect 8796 2728 10334 2736
rect 4824 2718 10334 2728
rect 2168 2714 10334 2718
rect -108 2662 10334 2714
rect -108 2654 9084 2662
rect -108 2644 5664 2654
rect 5718 2644 8172 2654
rect -108 2638 5658 2644
rect -108 2628 3732 2638
rect -108 2624 2840 2628
rect -108 2612 1888 2624
rect -108 2604 978 2612
rect -108 2532 142 2604
rect 242 2540 978 2604
rect 1078 2552 1888 2612
rect 1988 2552 2840 2624
rect 1078 2540 2840 2552
rect 242 2538 2840 2540
rect 2952 2548 3732 2628
rect 3844 2626 5658 2638
rect 3844 2548 4622 2626
rect 2952 2538 4622 2548
rect 242 2536 4622 2538
rect 4734 2542 5658 2626
rect 5764 2634 8172 2644
rect 5764 2542 6512 2634
rect 4734 2536 6512 2542
rect 242 2532 6512 2536
rect 6618 2532 7472 2634
rect 7578 2538 8172 2634
rect 8268 2546 9084 2654
rect 9180 2660 10334 2662
rect 9180 2546 10012 2660
rect 8268 2544 10012 2546
rect 10108 2544 10334 2660
rect 8268 2538 10334 2544
rect 7578 2532 10334 2538
rect -108 2470 10334 2532
rect -108 2468 2218 2470
rect 48 2344 166 2468
rect 48 2308 76 2344
rect 148 2308 166 2344
rect 48 2060 166 2308
rect 3582 2366 3688 2470
rect 4824 2468 10334 2470
rect 3582 2322 3596 2366
rect 3672 2322 3688 2366
rect 3582 2304 3688 2322
rect 6080 2330 6206 2468
rect 6080 2284 6100 2330
rect 6170 2284 6206 2330
rect 6080 2276 6206 2284
rect 2880 2264 4966 2272
rect 2880 2244 5688 2264
rect 2880 2210 2920 2244
rect 3288 2210 3378 2244
rect 3746 2210 3836 2244
rect 4204 2210 4294 2244
rect 4662 2236 5688 2244
rect 4662 2218 7540 2236
rect 4662 2210 5736 2218
rect 2880 2184 5736 2210
rect 6104 2184 6194 2218
rect 6562 2184 6652 2218
rect 7020 2184 7110 2218
rect 7478 2184 7540 2218
rect 2880 2178 7540 2184
rect 4858 2152 7540 2178
rect 8180 2080 8262 2468
rect 8786 2458 10334 2468
rect 8786 2352 8884 2458
rect 8786 2308 8800 2352
rect 8866 2308 8884 2352
rect 8786 2294 8884 2308
rect 2814 2062 4766 2076
rect 1438 2060 1728 2062
rect 48 2050 2002 2060
rect 48 1978 96 2050
rect 130 2046 2002 2050
rect 130 1978 1018 2046
rect 48 1974 1018 1978
rect 1052 1974 1932 2046
rect 1966 1974 2002 2046
rect 48 1972 2002 1974
rect 48 1964 1540 1972
rect 1624 1964 2002 1972
rect 2814 2052 2852 2062
rect 2888 2056 4766 2062
rect 2888 2052 3770 2056
rect 2814 1960 2844 2052
rect 2950 1974 3770 2052
rect 3806 1974 4684 2056
rect 4720 1974 4766 2056
rect 2950 1960 4766 1974
rect 2814 1946 4766 1960
rect 5634 2060 7596 2076
rect 5634 2056 7504 2060
rect 5634 2046 5672 2056
rect 5722 2052 7504 2056
rect 5634 1956 5662 2046
rect 5722 1966 6592 2052
rect 6632 1974 7504 2052
rect 7544 1974 7596 2060
rect 6632 1966 7596 1974
rect 5722 1964 7596 1966
rect 5716 1956 7596 1964
rect 5634 1944 7596 1956
rect 8176 2068 10088 2080
rect 8176 2058 10032 2068
rect 8176 2030 9124 2058
rect 8176 1968 8202 2030
rect 8238 1968 9124 2030
rect 8176 1966 9124 1968
rect 9162 1976 10032 2058
rect 10070 1976 10088 2068
rect 9162 1966 10088 1976
rect 8176 1928 10088 1966
rect 3296 1852 4288 1858
rect 3270 1844 4288 1852
rect 504 1742 1540 1764
rect 504 1736 1470 1742
rect 504 1664 560 1736
rect 594 1664 1470 1736
rect 1506 1664 1540 1742
rect 504 1642 1540 1664
rect 3270 1762 3310 1844
rect 3346 1838 4288 1844
rect 3346 1762 4238 1838
rect 3270 1756 4238 1762
rect 4274 1756 4288 1838
rect 3270 1724 4288 1756
rect 6102 1764 7128 1792
rect 1402 136 1534 1642
rect 98 119 1952 136
rect 98 85 159 119
rect 527 85 617 119
rect 985 85 1075 119
rect 1443 85 1533 119
rect 1901 85 1952 119
rect 98 48 1952 85
rect 1402 -132 1534 48
rect 3270 -132 3400 1724
rect 6102 1678 6134 1764
rect 6174 1678 7050 1764
rect 7090 1678 7128 1764
rect 8616 1718 9646 1722
rect 6102 1660 7128 1678
rect 8606 1686 9646 1718
rect 8606 1678 9558 1686
rect 6992 -128 7124 1660
rect 8606 1572 8636 1678
rect 8704 1580 9558 1678
rect 9626 1580 9646 1686
rect 8704 1572 9646 1580
rect 8606 1542 9646 1572
rect 8606 136 8728 1542
rect 8212 112 10048 136
rect 8212 78 8260 112
rect 8628 78 8718 112
rect 9086 78 9176 112
rect 9544 78 9634 112
rect 10002 78 10048 112
rect 8212 60 10048 78
rect 8606 -72 8728 60
rect 8606 -128 8726 -72
rect 1402 -164 3400 -132
rect 1402 -262 3406 -164
rect 6988 -212 8726 -128
rect 2302 -912 2520 -262
rect 1330 -1016 1404 -946
rect 2302 -948 2328 -912
rect 2468 -948 2520 -912
rect 2302 -962 2520 -948
rect 7798 -900 7912 -212
rect 7798 -940 7816 -900
rect 7900 -940 7912 -900
rect 7798 -954 7912 -940
rect 2298 -1008 2542 -992
rect 2298 -1054 2362 -1008
rect 2468 -1054 2542 -1008
rect 2298 -1116 2542 -1054
rect 2298 -1162 2354 -1116
rect 2460 -1162 2542 -1116
rect 2298 -1272 2542 -1162
rect 7790 -996 7926 -986
rect 7790 -1036 7816 -996
rect 7896 -1036 7926 -996
rect 8894 -1010 8962 -934
rect 7790 -1102 7926 -1036
rect 7790 -1142 7818 -1102
rect 7898 -1142 7926 -1102
rect 7790 -1272 7926 -1142
rect 2298 -1452 7940 -1272
rect 2298 -1458 2542 -1452
rect 5566 -2066 5858 -1452
rect 3710 -2072 8418 -2066
rect 3710 -2080 6508 -2072
rect 3710 -2084 5600 -2080
rect 3710 -2180 3766 -2084
rect 3814 -2092 5600 -2084
rect 3814 -2180 4682 -2092
rect 3710 -2188 4682 -2180
rect 4730 -2176 5600 -2092
rect 5648 -2168 6508 -2080
rect 6556 -2078 8418 -2072
rect 6556 -2168 7414 -2078
rect 5648 -2174 7414 -2168
rect 7462 -2174 8346 -2078
rect 8394 -2174 8418 -2078
rect 5648 -2176 8418 -2174
rect 4730 -2188 8418 -2176
rect 3710 -2198 8418 -2188
rect 5566 -2208 5858 -2198
rect 4146 -2256 8900 -2250
rect 4146 -2262 8784 -2256
rect 4146 -2274 6040 -2262
rect 4146 -2286 5122 -2274
rect 4146 -2396 4198 -2286
rect 4268 -2384 5122 -2286
rect 5192 -2284 6040 -2274
rect 6110 -2284 6964 -2262
rect 5192 -2384 6028 -2284
rect 6142 -2372 6964 -2284
rect 7034 -2274 8784 -2262
rect 7034 -2372 7888 -2274
rect 4268 -2392 6028 -2384
rect 6142 -2384 7888 -2372
rect 7958 -2366 8784 -2274
rect 8854 -2366 8900 -2256
rect 7958 -2384 8900 -2366
rect 6142 -2392 8900 -2384
rect 4268 -2396 8900 -2392
rect 4146 -2414 8900 -2396
rect 3328 -4427 8872 -4396
rect 3328 -4461 3835 -4427
rect 4203 -4461 4293 -4427
rect 4661 -4461 4751 -4427
rect 5119 -4461 5209 -4427
rect 5577 -4461 5667 -4427
rect 6035 -4461 6125 -4427
rect 6493 -4461 6583 -4427
rect 6951 -4461 7041 -4427
rect 7409 -4461 7499 -4427
rect 7867 -4461 7957 -4427
rect 8325 -4461 8415 -4427
rect 8783 -4461 8872 -4427
rect 3328 -4476 8872 -4461
rect 3328 -4480 3890 -4476
rect 7666 -4538 7842 -4510
rect 7666 -4572 7688 -4538
rect 7790 -4572 7842 -4538
rect 7666 -4692 7842 -4572
rect 3504 -4764 9152 -4692
rect 3504 -4770 6492 -4764
rect 3504 -4878 3716 -4770
rect 3830 -4786 5552 -4770
rect 3830 -4878 4662 -4786
rect 3504 -4894 4662 -4878
rect 4776 -4878 5552 -4786
rect 5666 -4788 6492 -4770
rect 5666 -4878 6028 -4788
rect 4776 -4894 6028 -4878
rect 3504 -4896 6028 -4894
rect 6142 -4872 6492 -4788
rect 6606 -4770 8314 -4764
rect 6606 -4872 7420 -4770
rect 6142 -4878 7420 -4872
rect 7534 -4872 8314 -4770
rect 8428 -4872 9152 -4764
rect 7534 -4878 9152 -4872
rect 6142 -4896 9152 -4878
rect 3504 -5042 9152 -4896
<< via1 >>
rect 5664 2644 5718 2654
rect 2840 2538 2952 2628
rect 5664 2564 5718 2644
rect 2844 1980 2852 2052
rect 2852 1980 2888 2052
rect 2888 1980 2950 2052
rect 2844 1960 2950 1980
rect 5662 1964 5672 2046
rect 5672 1964 5716 2046
rect 5662 1956 5716 1964
rect 6028 -2372 6040 -2284
rect 6040 -2372 6110 -2284
rect 6110 -2372 6142 -2284
rect 6028 -2392 6142 -2372
rect 6028 -4896 6142 -4788
<< metal2 >>
rect 2818 2628 2990 2722
rect 2818 2538 2840 2628
rect 2952 2538 2990 2628
rect 2818 2052 2990 2538
rect 2818 1960 2844 2052
rect 2950 1960 2990 2052
rect 2818 1920 2990 1960
rect 5648 2654 5734 2730
rect 5648 2564 5664 2654
rect 5718 2564 5734 2654
rect 5648 2046 5734 2564
rect 5648 1956 5662 2046
rect 5716 1956 5734 2046
rect 5648 1924 5734 1956
rect 6006 -2284 6188 -2262
rect 6006 -2392 6028 -2284
rect 6142 -2392 6188 -2284
rect 6006 -4788 6188 -2392
rect 6006 -4896 6028 -4788
rect 6142 -4896 6188 -4788
rect 6006 -4904 6188 -4896
use sky130_fd_pr__nfet_01v8_lvt_V62P9P  sky130_fd_pr__nfet_01v8_lvt_V62P9P_0
timestamp 1606420870
transform 1 0 6309 0 1 -3189
box -2686 -1410 2686 1410
use sky130_fd_pr__nfet_01v8_lvt_6NXDEK  sky130_fd_pr__nfet_01v8_lvt_6NXDEK_1
timestamp 1606420870
transform 0 1 7874 -1 0 -971
box -211 -1210 211 1210
use sky130_fd_pr__nfet_01v8_lvt_6NXDEK  sky130_fd_pr__nfet_01v8_lvt_6NXDEK_0
timestamp 1606420870
transform 0 1 2424 -1 0 -981
box -211 -1210 211 1210
use sky130_fd_pr__pfet_01v8_lvt_AG2VEQ  sky130_fd_pr__pfet_01v8_lvt_AG2VEQ_2
timestamp 1606420870
transform 1 0 9131 0 1 1159
box -1083 -1219 1083 1219
use sky130_fd_pr__pfet_01v8_lvt_AG2VEQ  sky130_fd_pr__pfet_01v8_lvt_AG2VEQ_1
timestamp 1606420870
transform 1 0 6607 0 1 1137
box -1083 -1219 1083 1219
use sky130_fd_pr__pfet_01v8_AG284Q  sky130_fd_pr__pfet_01v8_AG284Q_0
timestamp 1606420870
transform 1 0 3791 0 1 1163
box -1083 -1219 1083 1219
use sky130_fd_pr__pfet_01v8_lvt_AG2VEQ  sky130_fd_pr__pfet_01v8_lvt_AG2VEQ_0
timestamp 1606420870
transform 1 0 1037 0 1 1169
box -1083 -1219 1083 1219
<< labels >>
rlabel metal1 1118 2480 1338 2708 1 Vdd
port 1 n
rlabel metal1 1456 -132 1528 -70 1 D2l
port 2 n
rlabel metal1 5194 2196 5324 2246 1 Vctrl
port 3 n
rlabel metal1 2316 -232 2506 -150 1 D1l
port 4 n
rlabel metal1 7808 -204 7896 -136 1 D1r
port 5 n
rlabel metal1 1336 -1006 1394 -950 1 inp
port 6 n
rlabel metal1 8900 -998 8954 -952 1 inn
port 7 n
rlabel metal1 3346 -4468 3438 -4398 1 vbn
port 8 n
rlabel metal1 5802 -4912 5960 -4796 1 Gnd
port 9 n
<< end >>
