magic
tech sky130A
magscale 1 2
timestamp 1606359646
<< locali >>
rect 3174 662 3226 664
rect -102 618 3226 662
rect -102 614 3132 618
rect -100 366 -52 614
rect -100 332 28 366
rect 440 216 612 260
rect 740 254 954 260
rect 754 220 954 254
rect 1092 252 1308 260
rect 740 218 954 220
rect 1102 218 1308 252
rect 1446 252 1662 260
rect 1448 218 1662 252
rect 1092 216 1308 218
rect 1446 216 1662 218
rect 1796 216 2012 260
rect 2148 254 2364 260
rect 2500 254 2716 260
rect 3174 258 3226 618
rect 2150 220 2364 254
rect 2148 216 2364 220
rect 2504 220 2716 254
rect 2500 216 2716 220
rect 2852 220 3226 258
rect 2852 216 3180 220
<< viali >>
rect 32 340 66 374
rect 202 218 242 254
rect 402 216 436 250
rect 616 215 650 249
rect 720 220 754 254
rect 962 220 996 254
rect 1068 218 1102 252
rect 1314 222 1348 256
rect 1414 218 1448 252
rect 1664 220 1698 254
rect 1762 220 1796 254
rect 2016 220 2050 254
rect 2116 220 2150 254
rect 2376 218 2410 252
rect 2470 220 2504 254
rect 2728 215 2762 249
rect 2818 216 2852 250
<< metal1 >>
rect 3172 708 3272 714
rect -100 672 3272 708
rect -106 622 3272 672
rect -106 390 -36 622
rect 4 498 1630 594
rect 1634 496 3118 592
rect -106 374 86 390
rect -106 340 32 374
rect 66 340 86 374
rect -106 324 86 340
rect -112 254 256 260
rect -112 218 202 254
rect 242 218 256 254
rect -112 212 256 218
rect 390 250 666 262
rect 390 216 402 250
rect 436 249 666 250
rect 436 216 616 249
rect 390 215 616 216
rect 650 215 666 249
rect 390 200 666 215
rect 698 254 1020 266
rect 698 220 720 254
rect 754 220 962 254
rect 996 220 1020 254
rect 698 198 1020 220
rect 1052 256 1372 264
rect 1052 252 1314 256
rect 1052 218 1068 252
rect 1102 222 1314 252
rect 1348 222 1372 256
rect 1102 218 1372 222
rect 1052 196 1372 218
rect 1400 254 1720 266
rect 1400 252 1664 254
rect 1400 218 1414 252
rect 1448 220 1664 252
rect 1698 220 1720 254
rect 1448 218 1720 220
rect 1400 198 1720 218
rect 1756 254 2076 266
rect 1756 220 1762 254
rect 1796 220 2016 254
rect 2050 220 2076 254
rect 1756 198 2076 220
rect 2106 254 2426 268
rect 2106 220 2116 254
rect 2150 252 2426 254
rect 2150 220 2376 252
rect 2106 218 2376 220
rect 2410 218 2426 252
rect 2106 200 2426 218
rect 2462 254 2782 268
rect 3172 264 3272 622
rect 2462 220 2470 254
rect 2504 249 2782 254
rect 2504 220 2728 249
rect 2462 215 2728 220
rect 2762 215 2782 249
rect 2462 200 2782 215
rect 2812 250 3272 264
rect 2812 216 2818 250
rect 2852 216 3272 250
rect 2812 188 3272 216
rect 2 -48 3118 48
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1606359646
transform 1 0 2648 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1606359646
transform 1 0 2296 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1606359646
transform 1 0 1944 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1606359646
transform 1 0 1592 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1606359646
transform 1 0 1240 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1606359646
transform 1 0 888 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1606359646
transform 1 0 536 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1606359646
transform 1 0 3000 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0
timestamp 1606359646
transform 1 0 0 0 1 0
box -38 -48 498 592
<< labels >>
rlabel metal1 -96 226 -90 230 1 en
port 3 n
rlabel metal1 480 536 486 540 1 Vdd
port 1 n
rlabel metal1 480 -4 486 0 1 Gnd
port 2 n
rlabel metal1 -84 342 -70 362 1 out
port 4 n
<< end >>
