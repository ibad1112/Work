magic
tech sky130A
magscale 1 2
timestamp 1606076054
<< nwell >>
rect 5184 2660 5398 2676
rect -152 2404 5398 2660
rect -152 2384 5370 2404
<< nsubdiff >>
rect -84 2576 5344 2612
rect -84 2484 184 2576
rect 268 2572 1198 2576
rect 268 2484 492 2572
rect -84 2480 492 2484
rect 576 2480 834 2572
rect 918 2484 1198 2572
rect 1282 2572 1928 2576
rect 1282 2484 1550 2572
rect 918 2480 1550 2484
rect 1634 2484 1928 2572
rect 2012 2572 2622 2576
rect 2012 2484 2248 2572
rect 1634 2480 2248 2484
rect 2332 2484 2622 2572
rect 2706 2484 2968 2576
rect 3052 2572 4836 2576
rect 3052 2566 4346 2572
rect 3052 2484 3684 2566
rect 2332 2480 3684 2484
rect -84 2474 3684 2480
rect 3768 2480 4346 2566
rect 4430 2484 4836 2572
rect 4920 2484 5344 2576
rect 4430 2480 5344 2484
rect 3768 2474 5344 2480
rect -84 2452 5344 2474
<< nsubdiffcont >>
rect 184 2484 268 2576
rect 492 2480 576 2572
rect 834 2480 918 2572
rect 1198 2484 1282 2576
rect 1550 2480 1634 2572
rect 1928 2484 2012 2576
rect 2248 2480 2332 2572
rect 2622 2484 2706 2576
rect 2968 2484 3052 2576
rect 3684 2474 3768 2566
rect 4346 2480 4430 2572
rect 4836 2484 4920 2576
<< locali >>
rect -20 2564 184 2576
rect -20 2490 56 2564
rect 140 2490 184 2564
rect -20 2484 184 2490
rect 268 2572 1198 2576
rect 268 2570 492 2572
rect 268 2496 344 2570
rect 428 2496 492 2570
rect 268 2484 492 2496
rect -20 2480 492 2484
rect 576 2570 834 2572
rect 576 2496 668 2570
rect 752 2496 834 2570
rect 576 2480 834 2496
rect 918 2570 1198 2572
rect 918 2496 1016 2570
rect 1100 2496 1198 2570
rect 918 2484 1198 2496
rect 1282 2574 1928 2576
rect 1282 2572 1746 2574
rect 1282 2570 1550 2572
rect 1282 2496 1390 2570
rect 1474 2496 1550 2570
rect 1282 2484 1550 2496
rect 918 2480 1550 2484
rect 1634 2500 1746 2572
rect 1830 2500 1928 2574
rect 1634 2484 1928 2500
rect 2012 2572 2622 2576
rect 2012 2564 2248 2572
rect 2012 2490 2062 2564
rect 2146 2490 2248 2564
rect 2012 2484 2248 2490
rect 1634 2480 2248 2484
rect 2332 2570 2622 2572
rect 2332 2496 2484 2570
rect 2568 2496 2622 2570
rect 2332 2484 2622 2496
rect 2706 2574 2968 2576
rect 2706 2500 2804 2574
rect 2888 2500 2968 2574
rect 2706 2484 2968 2500
rect 3052 2570 3882 2576
rect 3052 2496 3118 2570
rect 3202 2496 3470 2570
rect 3554 2566 3882 2570
rect 3554 2496 3684 2566
rect 3052 2484 3684 2496
rect 2332 2480 3684 2484
rect -20 2474 3684 2480
rect 3768 2506 3882 2566
rect 3966 2574 4836 2576
rect 3966 2572 4720 2574
rect 3966 2570 4346 2572
rect 3966 2506 4212 2570
rect 3768 2496 4212 2506
rect 4296 2496 4346 2570
rect 3768 2480 4346 2496
rect 4430 2570 4720 2572
rect 4430 2496 4452 2570
rect 4536 2500 4720 2570
rect 4804 2500 4836 2574
rect 4536 2496 4836 2500
rect 4430 2484 4836 2496
rect 4920 2570 5316 2576
rect 4920 2496 4944 2570
rect 5028 2496 5316 2570
rect 4920 2484 5316 2496
rect 4430 2480 5316 2484
rect 3768 2474 5316 2480
rect 1204 2470 3808 2474
rect 1204 2314 1264 2470
rect 3746 2322 3806 2470
rect 3270 2004 3304 2088
rect 3586 2012 3620 2096
rect 3902 2016 3936 2100
<< viali >>
rect 56 2490 140 2564
rect 344 2496 428 2570
rect 668 2496 752 2570
rect 1016 2496 1100 2570
rect 1390 2496 1474 2570
rect 1746 2500 1830 2574
rect 2062 2490 2146 2564
rect 2484 2496 2568 2570
rect 2804 2500 2888 2574
rect 3118 2496 3202 2570
rect 3470 2496 3554 2570
rect 3882 2506 3966 2580
rect 4212 2496 4296 2570
rect 4452 2496 4536 2570
rect 4720 2500 4804 2574
rect 4944 2496 5028 2570
rect 159 2213 227 2247
rect 317 2213 385 2247
rect 475 2213 543 2247
rect 633 2213 701 2247
rect 791 2213 859 2247
rect 949 2213 1017 2247
rect 1107 2213 1175 2247
rect 1265 2213 1333 2247
rect 1423 2213 1491 2247
rect 1581 2213 1649 2247
rect 1739 2213 1807 2247
rect 1897 2213 1965 2247
rect 2055 2213 2123 2247
rect 2213 2213 2281 2247
rect 2371 2213 2439 2247
rect 2860 2218 2928 2252
rect 3018 2218 3086 2252
rect 3176 2218 3244 2252
rect 3334 2218 3402 2252
rect 3492 2218 3560 2252
rect 3650 2218 3718 2252
rect 3808 2218 3876 2252
rect 3966 2218 4034 2252
rect 4124 2218 4192 2252
rect 4282 2218 4350 2252
rect 4440 2218 4508 2252
rect 4598 2218 4666 2252
rect 4756 2218 4824 2252
rect 4914 2218 4982 2252
rect 5072 2218 5140 2252
rect 98 2000 136 2070
rect 414 2008 452 2078
rect 726 2008 764 2078
rect 1044 2014 1082 2084
rect 1358 2006 1396 2076
rect 1676 2002 1714 2072
rect 1992 2008 2030 2078
rect 2308 2012 2346 2082
rect 2796 1958 2832 2060
rect 3110 1972 3146 2074
rect 3428 1972 3464 2074
rect 3746 1968 3782 2070
rect 4058 1974 4094 2076
rect 4374 1976 4410 2078
rect 4690 1968 4726 2070
rect 5012 1972 5048 2074
rect 252 1746 290 1816
rect 566 1750 604 1820
rect 888 1748 926 1818
rect 1204 1752 1242 1822
rect 1522 1756 1560 1826
rect 1834 1756 1872 1826
rect 2156 1756 2194 1826
rect 2466 1752 2504 1822
rect 2956 1742 2990 1850
rect 3268 1750 3302 1858
rect 3586 1746 3620 1854
rect 3902 1748 3936 1856
rect 4222 1748 4256 1856
rect 4536 1742 4570 1850
rect 4852 1742 4886 1850
rect 5168 1742 5202 1850
rect 2371 85 2439 119
rect 2392 -402 2452 -368
rect 2894 -404 2954 -370
rect 2392 -490 2452 -456
rect 2894 -492 2954 -458
rect 2396 -602 2462 -568
rect 2892 -606 2958 -572
rect 2642 -1016 2688 -982
rect 1478 -1586 1530 -1552
rect 1810 -1592 1862 -1558
rect 2292 -1592 2344 -1558
rect 2944 -1586 2996 -1552
rect 3530 -1590 3582 -1556
rect 3848 -1588 3900 -1554
<< metal1 >>
rect -110 2592 5338 2628
rect -110 2564 66 2592
rect 172 2580 5338 2592
rect 172 2574 3882 2580
rect 172 2570 1746 2574
rect -110 2490 56 2564
rect 172 2496 344 2570
rect 428 2496 668 2570
rect 752 2496 1016 2570
rect 1100 2496 1390 2570
rect 1474 2500 1746 2570
rect 1830 2570 2804 2574
rect 1830 2564 2484 2570
rect 1830 2500 2062 2564
rect 1474 2496 2062 2500
rect 172 2490 2062 2496
rect 2146 2496 2484 2564
rect 2568 2500 2804 2570
rect 2888 2570 3882 2574
rect 2888 2500 3118 2570
rect 2568 2496 3118 2500
rect 3202 2496 3470 2570
rect 3554 2506 3882 2570
rect 3966 2574 5338 2580
rect 3966 2570 4720 2574
rect 3966 2506 4212 2570
rect 3554 2496 4212 2506
rect 4296 2496 4452 2570
rect 4536 2500 4720 2570
rect 4804 2570 5338 2574
rect 4804 2500 4944 2570
rect 4536 2496 4944 2500
rect 5028 2566 5338 2570
rect 5028 2496 5132 2566
rect 2146 2490 5132 2496
rect -110 2458 66 2490
rect 172 2474 5132 2490
rect 5234 2474 5338 2566
rect 172 2458 5338 2474
rect -110 2436 5338 2458
rect 2830 2274 5170 2278
rect 132 2252 5170 2274
rect 132 2247 2860 2252
rect 132 2213 159 2247
rect 227 2213 317 2247
rect 385 2213 475 2247
rect 543 2213 633 2247
rect 701 2213 791 2247
rect 859 2213 949 2247
rect 1017 2213 1107 2247
rect 1175 2213 1265 2247
rect 1333 2213 1423 2247
rect 1491 2213 1581 2247
rect 1649 2213 1739 2247
rect 1807 2213 1897 2247
rect 1965 2213 2055 2247
rect 2123 2213 2213 2247
rect 2281 2213 2371 2247
rect 2439 2218 2860 2247
rect 2928 2218 3018 2252
rect 3086 2218 3176 2252
rect 3244 2218 3334 2252
rect 3402 2218 3492 2252
rect 3560 2218 3650 2252
rect 3718 2218 3808 2252
rect 3876 2218 3966 2252
rect 4034 2218 4124 2252
rect 4192 2218 4282 2252
rect 4350 2218 4440 2252
rect 4508 2218 4598 2252
rect 4666 2218 4756 2252
rect 4824 2218 4914 2252
rect 4982 2218 5072 2252
rect 5140 2218 5170 2252
rect 2439 2213 5170 2218
rect 132 2200 5170 2213
rect 2350 2196 3320 2200
rect 26 2112 234 2124
rect 26 1978 66 2112
rect 172 2110 234 2112
rect 172 2084 2356 2110
rect 172 2078 1044 2084
rect 172 2008 414 2078
rect 452 2008 726 2078
rect 764 2014 1044 2078
rect 1082 2082 2356 2084
rect 1082 2078 2308 2082
rect 1082 2076 1992 2078
rect 1082 2014 1358 2076
rect 764 2008 1358 2014
rect 172 2006 1358 2008
rect 1396 2072 1992 2076
rect 1396 2006 1676 2072
rect 172 2002 1676 2006
rect 1714 2008 1992 2072
rect 2030 2012 2308 2078
rect 2346 2012 2356 2082
rect 2030 2008 2356 2012
rect 1714 2002 2356 2008
rect 172 1978 2356 2002
rect 26 1962 2356 1978
rect 26 1944 234 1962
rect 2750 2084 2874 2086
rect 2750 2078 5062 2084
rect 2750 2076 4374 2078
rect 2750 2074 4058 2076
rect 2750 2060 3110 2074
rect 2750 1958 2796 2060
rect 2832 1972 3110 2060
rect 3146 1972 3428 2074
rect 3464 2070 4058 2074
rect 3464 1972 3746 2070
rect 2832 1968 3746 1972
rect 3782 1974 4058 2070
rect 4094 1976 4374 2076
rect 4410 2074 5062 2078
rect 4410 2070 5012 2074
rect 4410 1976 4690 2070
rect 4094 1974 4690 1976
rect 3782 1968 4690 1974
rect 4726 1972 5012 2070
rect 5048 1972 5062 2074
rect 4726 1968 5062 1972
rect 2832 1958 5062 1968
rect 2750 1950 5062 1958
rect 2426 1864 2546 1870
rect 238 1826 2546 1864
rect 2750 1832 2874 1950
rect 5108 1864 5260 1878
rect 238 1822 1522 1826
rect 238 1820 1204 1822
rect 238 1816 566 1820
rect 238 1746 252 1816
rect 290 1750 566 1816
rect 604 1818 1204 1820
rect 604 1750 888 1818
rect 290 1748 888 1750
rect 926 1752 1204 1818
rect 1242 1756 1522 1822
rect 1560 1756 1834 1826
rect 1872 1756 2156 1826
rect 2194 1822 2546 1826
rect 2194 1756 2466 1822
rect 1242 1752 2466 1756
rect 2504 1752 2546 1822
rect 926 1748 2546 1752
rect 290 1746 2546 1748
rect 238 1700 2546 1746
rect 2426 134 2546 1700
rect 2352 119 2546 134
rect 2352 85 2371 119
rect 2439 85 2546 119
rect 2352 64 2546 85
rect 2426 -152 2546 64
rect 2372 -178 2546 -152
rect 2738 62 2874 1832
rect 2944 1858 5260 1864
rect 2944 1850 3268 1858
rect 2944 1742 2956 1850
rect 2990 1750 3268 1850
rect 3302 1856 5260 1858
rect 3302 1854 3902 1856
rect 3302 1750 3586 1854
rect 2990 1746 3586 1750
rect 3620 1748 3902 1854
rect 3936 1748 4222 1856
rect 4256 1850 5260 1856
rect 4256 1748 4536 1850
rect 3620 1746 4536 1748
rect 2990 1742 4536 1746
rect 4570 1742 4852 1850
rect 4886 1840 5168 1850
rect 5202 1840 5260 1850
rect 4886 1748 5150 1840
rect 5252 1748 5260 1840
rect 4886 1742 5168 1748
rect 5202 1742 5260 1748
rect 2944 1734 5260 1742
rect 5108 1724 5260 1734
rect 2738 -136 2862 62
rect 2372 -352 2474 -178
rect 2738 -192 2976 -136
rect 2846 -196 2976 -192
rect 2372 -368 2478 -352
rect 2372 -402 2392 -368
rect 2452 -402 2478 -368
rect 2372 -406 2478 -402
rect 2378 -410 2478 -406
rect 2874 -370 2976 -196
rect 2874 -404 2894 -370
rect 2954 -404 2976 -370
rect 2874 -410 2976 -404
rect 2366 -456 2476 -450
rect 2366 -490 2392 -456
rect 2452 -490 2476 -456
rect 2366 -558 2476 -490
rect 2872 -458 2982 -452
rect 2872 -492 2894 -458
rect 2954 -492 2982 -458
rect 2872 -558 2982 -492
rect 2362 -568 2982 -558
rect 2362 -602 2396 -568
rect 2462 -572 2982 -568
rect 2462 -602 2892 -572
rect 2362 -606 2892 -602
rect 2958 -606 2982 -572
rect 2362 -620 2982 -606
rect 2622 -728 2708 -620
rect 2622 -982 2706 -728
rect 2622 -1016 2642 -982
rect 2688 -1016 2706 -982
rect 2622 -1018 2706 -1016
rect 2626 -1022 2706 -1018
rect 1170 -1552 4300 -1522
rect 1170 -1586 1478 -1552
rect 1530 -1558 2944 -1552
rect 1530 -1586 1810 -1558
rect 1170 -1592 1810 -1586
rect 1862 -1592 2292 -1558
rect 2344 -1586 2944 -1558
rect 2996 -1554 4300 -1552
rect 2996 -1556 3848 -1554
rect 2996 -1586 3530 -1556
rect 2344 -1590 3530 -1586
rect 3582 -1588 3848 -1556
rect 3900 -1588 4300 -1554
rect 3582 -1590 4300 -1588
rect 2344 -1592 4300 -1590
rect 1170 -1748 4300 -1592
<< rmetal1 >>
rect 234 1960 2356 1962
<< via1 >>
rect 66 2564 172 2592
rect 66 2490 140 2564
rect 140 2490 172 2564
rect 66 2458 172 2490
rect 5132 2474 5234 2566
rect 66 2070 172 2112
rect 66 2000 98 2070
rect 98 2000 136 2070
rect 136 2000 172 2070
rect 66 1978 172 2000
rect 5150 1748 5168 1840
rect 5168 1748 5202 1840
rect 5202 1748 5252 1840
<< metal2 >>
rect 44 2592 194 2618
rect 44 2458 66 2592
rect 172 2458 194 2592
rect 44 2112 194 2458
rect 44 1978 66 2112
rect 172 1978 194 2112
rect 44 1938 194 1978
rect 5116 2566 5276 2584
rect 5116 2474 5132 2566
rect 5234 2474 5276 2566
rect 5116 1840 5276 2474
rect 5116 1748 5150 1840
rect 5252 1748 5276 1840
rect 5116 1724 5276 1748
use sky130_fd_pr__pfet_01v8_NC6LGM  sky130_fd_pr__pfet_01v8_NC6LGM_0
timestamp 1606057846
transform 1 0 1299 0 1 1166
box -1352 -1219 1352 1219
use sky130_fd_pr__pfet_01v8_NC6LGM  sky130_fd_pr__pfet_01v8_NC6LGM_1
timestamp 1606057846
transform 1 0 4000 0 1 1171
box -1352 -1219 1352 1219
use sky130_fd_pr__nfet_01v8_lvt_D42ZUM  sky130_fd_pr__nfet_01v8_lvt_D42ZUM_0
timestamp 1606076054
transform 0 1 2924 -1 0 -431
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_D42ZUM  sky130_fd_pr__nfet_01v8_lvt_D42ZUM_1
timestamp 1606076054
transform 0 1 2422 -1 0 -429
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_69NU8X  sky130_fd_pr__nfet_01v8_lvt_69NU8X_0
timestamp 1606076054
transform 0 1 2704 -1 0 -1228
box -396 -1470 396 1470
<< labels >>
rlabel metal1 2356 2494 2412 2550 1 Vdd
port 1 n
rlabel metal1 2460 -134 2516 -78 1 ON2b
port 2 n
rlabel metal1 2778 -132 2834 -76 1 ON1b
port 3 n
rlabel space 2314 -438 2330 -418 1 ON1a
port 4 n
rlabel space 3010 -442 3026 -422 1 ON2a
port 5 n
rlabel metal1 2664 -1694 2750 -1640 1 Gnd
port 6 n
rlabel metal1 2652 -744 2684 -700 1 Itail_b
rlabel space 1370 -1286 1410 -1216 1 vbiasn
port 7 n
<< end >>
